Group|Creator|Element|VR|VM|Name
0019|1.2.840.113681|10|ST|1|CRImageParamsCommon
0019|1.2.840.113681|11|ST|1|CRImageIPParamsSingle
0019|1.2.840.113681|12|ST|1|CRImageIPParamsLeft
0019|1.2.840.113681|13|ST|1|CRImageIPParamsRight
0087|1.2.840.113708.794.1.1.2.0|10|CS|1|MediaType
0087|1.2.840.113708.794.1.1.2.0|20|CS|1|MediaLocation
0087|1.2.840.113708.794.1.1.2.0|50|IS|1|EstimatedRetrieveTime
0009|ACUSON|00|IS|1|Unknown
0009|ACUSON|01|IS|1|Unknown
0009|ACUSON|02|UN|1|Unknown
0009|ACUSON|03|UN|1|Unknown
0009|ACUSON|04|UN|1|Unknown
0009|ACUSON|05|UN|1|Unknown
0009|ACUSON|06|UN|1|Unknown
0009|ACUSON|07|UN|1|Unknown
0009|ACUSON|08|LT|1|Unknown
0009|ACUSON|09|LT|1|Unknown
0009|ACUSON|0a|IS|1|Unknown
0009|ACUSON|0b|IS|1|Unknown
0009|ACUSON|0c|IS|1|Unknown
0009|ACUSON|0d|IS|1|Unknown
0009|ACUSON|0e|IS|1|Unknown
0009|ACUSON|0f|UN|1|Unknown
0009|ACUSON|10|IS|1|Unknown
0009|ACUSON|11|UN|1|Unknown
0009|ACUSON|12|IS|1|Unknown
0009|ACUSON|13|IS|1|Unknown
0009|ACUSON|14|LT|1|Unknown
0009|ACUSON|15|UN|1|Unknown
0003|AEGIS_DICOM_2.00|00|US|1-n|Unknown
0005|AEGIS_DICOM_2.00|00|US|1-n|Unknown
0009|AEGIS_DICOM_2.00|00|US|1-n|Unknown
0019|AEGIS_DICOM_2.00|00|US|1-n|Unknown
0029|AEGIS_DICOM_2.00|00|US|1-n|Unknown
1369|AEGIS_DICOM_2.00|00|US|1-n|Unknown
0009|AGFA|10|LO|1|Unknown
0009|AGFA|11|LO|1|Unknown
0009|AGFA|13|LO|1|Unknown
0009|AGFA|14|LO|1|Unknown
0009|AGFA|15|LO|1|Unknown
0029|CAMTRONICS IP|10|LT|1|Unknown
0029|CAMTRONICS IP|20|UN|1|Unknown
0029|CAMTRONICS IP|30|UN|1|Unknown
0029|CAMTRONICS IP|40|UN|1|Unknown
0029|CAMTRONICS|10|LT|1|Commentline
0029|CAMTRONICS|20|DS|1|EdgeEnhancementCoefficient
0029|CAMTRONICS|50|LT|1|SceneText
0029|CAMTRONICS|60|LT|1|ImageText
0029|CAMTRONICS|70|IS|1|PixelShiftHorizontal
0029|CAMTRONICS|80|IS|1|PixelShiftVertical
0029|CAMTRONICS|90|IS|1|Unknown
0009|CARDIO-D.R. 1.0|00|UL|1|FileLocation
0009|CARDIO-D.R. 1.0|01|UL|1|FileSize
0009|CARDIO-D.R. 1.0|40|SQ|1|AlternateImageSequence
0019|CARDIO-D.R. 1.0|00|CS|1|ImageBlankingShape
0019|CARDIO-D.R. 1.0|02|IS|1|ImageBlankingLeftVerticalEdge
0019|CARDIO-D.R. 1.0|04|IS|1|ImageBlankingRightVerticalEdge
0019|CARDIO-D.R. 1.0|06|IS|1|ImageBlankingUpperHorizontalEdge
0019|CARDIO-D.R. 1.0|08|IS|1|ImageBlankingLowerHorizontalEdge
0019|CARDIO-D.R. 1.0|10|IS|1|CenterOfCircularImageBlanking
0019|CARDIO-D.R. 1.0|12|IS|1|RadiusOfCircularImageBlanking
0019|CARDIO-D.R. 1.0|30|UL|1|MaximumImageFrameSize
0021|CARDIO-D.R. 1.0|13|IS|1|ImageSequenceNumber
0119|MRSC|1502|TM|1|SERTime
0029|CARDIO-D.R. 1.0|00|SQ|1|EdgeEnhancementSequence
0029|CARDIO-D.R. 1.0|01|US|2|ConvolutionKernelSize
0029|CARDIO-D.R. 1.0|02|DS|1-n|ConvolutionKernelCoefficients
0029|CARDIO-D.R. 1.0|03|DS|1|EdgeEnhancementGain
0025|CMR42 CIRCLECVI|1010|LO|1|WorkspaceID
0025|CMR42 CIRCLECVI|1020|LO|1|WorkspaceTimeString
0025|CMR42 CIRCLECVI|1030|OB|1|WorkspaceStream
0009|DCMTK_ANONYMIZER|00|SQ|1|AnonymizerUIDMap
0009|DCMTK_ANONYMIZER|10|UI|1|AnonymizerUIDKey
0009|DCMTK_ANONYMIZER|20|UI|1|AnonymizerUIDValue
0009|DCMTK_ANONYMIZER|30|SQ|1|AnonymizerPatientIDMap
0009|DCMTK_ANONYMIZER|40|LO|1|AnonymizerPatientIDKey
0009|DCMTK_ANONYMIZER|50|LO|1|AnonymizerPatientIDValue
0019|DIDI TO PCR 1.1|22|UN|1|RouteAET
0019|DIDI TO PCR 1.1|23|DS|1|PCRPrintScale
0019|DIDI TO PCR 1.1|24|UN|1|PCRPrintJobEnd
0019|DIDI TO PCR 1.1|25|IS|1|PCRNoFilmCopies
0019|DIDI TO PCR 1.1|26|IS|1|PCRFilmLayoutPosition
0019|DIDI TO PCR 1.1|27|UN|1|PCRPrintReportName
0019|DIDI TO PCR 1.1|70|UN|1|RADProtocolPrinter
0019|DIDI TO PCR 1.1|71|UN|1|RADProtocolMedium
0019|DIDI TO PCR 1.1|90|LO|1|UnprocessedFlag
0019|DIDI TO PCR 1.1|91|UN|1|KeyValues
0019|DIDI TO PCR 1.1|92|UN|1|DestinationPostprocessingFunction
0019|DIDI TO PCR 1.1|A0|UN|1|Version
0019|DIDI TO PCR 1.1|A1|UN|1|RangingMode
0019|DIDI TO PCR 1.1|A2|UN|1|AbdomenBrightness
0019|DIDI TO PCR 1.1|A3|UN|1|FixedBrightness
0019|DIDI TO PCR 1.1|A4|UN|1|DetailContrast
0019|DIDI TO PCR 1.1|A5|UN|1|ContrastBalance
0019|DIDI TO PCR 1.1|A6|UN|1|StructureBoost
0019|DIDI TO PCR 1.1|A7|UN|1|StructurePreference
0019|DIDI TO PCR 1.1|A8|UN|1|NoiseRobustness
0019|DIDI TO PCR 1.1|A9|UN|1|NoiseDoseLimit
0019|DIDI TO PCR 1.1|AA|UN|1|NoiseDoseStep
0019|DIDI TO PCR 1.1|AB|UN|1|NoiseFrequencyLimit
0019|DIDI TO PCR 1.1|AC|UN|1|WeakContrastLimit
0019|DIDI TO PCR 1.1|AD|UN|1|StrongContrastLimit
0019|DIDI TO PCR 1.1|AE|UN|1|StructureBoostOffset
0019|DIDI TO PCR 1.1|AF|UN|1|SmoothGain
0019|DIDI TO PCR 1.1|B0|UN|1|MeasureField1
0019|DIDI TO PCR 1.1|B1|UN|1|MeasureField2
0019|DIDI TO PCR 1.1|B2|UN|1|KeyPercentile1
0019|DIDI TO PCR 1.1|B3|UN|1|KeyPercentile2
0019|DIDI TO PCR 1.1|B4|UN|1|DensityLUT
0019|DIDI TO PCR 1.1|B5|UN|1|Brightness
0019|DIDI TO PCR 1.1|B6|UN|1|Gamma
0089|DIDI TO PCR 1.1|10|SQ|1|Unknown
0029|DIGISCAN IMAGE|31|US|1-n|Unknown
0029|DIGISCAN IMAGE|32|US|1-n|Unknown
0029|DIGISCAN IMAGE|33|LT|1|Unknown
0029|DIGISCAN IMAGE|34|LT|1|Unknown
0015|DLX_EXAMS_01|01|DS|1|StenosisCalibrationRatio
0015|DLX_EXAMS_01|02|DS|1|StenosisMagnification
0015|DLX_EXAMS_01|03|DS|1|CardiacCalibrationRatio
0011|DLX_PATNT_01|01|LT|1|PatientDOB
0019|DLX_SERIE_01|01|DS|1|AngleValueLArm
0019|DLX_SERIE_01|02|DS|1|AngleValuePArm
0019|DLX_SERIE_01|03|DS|1|AngleValueCArm
0019|DLX_SERIE_01|04|CS|1|AngleLabelLArm
0019|DLX_SERIE_01|05|CS|1|AngleLabelPArm
0019|DLX_SERIE_01|06|CS|1|AngleLabelCArm
0019|DLX_SERIE_01|07|ST|1|ProcedureName
0019|DLX_SERIE_01|08|ST|1|ExamName
0019|DLX_SERIE_01|09|SH|1|PatientSize
0019|DLX_SERIE_01|0a|IS|1|RecordView
0019|DLX_SERIE_01|10|DS|1|InjectorDelay
0019|DLX_SERIE_01|11|CS|1|AutoInject
0019|DLX_SERIE_01|14|IS|1|AcquisitionMode
0019|DLX_SERIE_01|15|CS|1|CameraRotationEnabled
0019|DLX_SERIE_01|16|CS|1|ReverseSweep
0019|DLX_SERIE_01|17|IS|1|SpatialFilterStrength
0019|DLX_SERIE_01|18|IS|1|ZoomFactor
0019|DLX_SERIE_01|19|IS|1|XZoomCenter
0019|DLX_SERIE_01|1a|IS|1|YZoomCenter
0019|DLX_SERIE_01|1b|DS|1|Focus
0019|DLX_SERIE_01|1c|CS|1|Dose
0019|DLX_SERIE_01|1d|IS|1|SideMark
0019|DLX_SERIE_01|1e|IS|1|PercentageLandscape
0019|DLX_SERIE_01|1f|DS|1|ExposureDuration
00E1|ELSCINT1|01|US|1|DataDictionaryVersion
00E1|ELSCINT1|14|LT|1|Unknown
00E1|ELSCINT1|22|DS|2|Unknown
00E1|ELSCINT1|23|DS|2|Unknown
00E1|ELSCINT1|24|LT|1|Unknown
00E1|ELSCINT1|25|LT|1|Unknown
00E1|ELSCINT1|40|SH|1|OffsetFromCTMRImages
0601|ELSCINT1|00|SH|1|ImplementationVersion
0601|ELSCINT1|20|DS|1|RelativeTablePosition
0601|ELSCINT1|21|DS|1|RelativeTableHeight
0601|ELSCINT1|30|SH|1|SurviewDirection
0601|ELSCINT1|31|DS|1|SurviewLength
0601|ELSCINT1|50|SH|1|ImageViewType
0601|ELSCINT1|70|DS|1|BatchNumber
0601|ELSCINT1|71|DS|1|BatchSize
0601|ELSCINT1|72|DS|1|BatchSliceNumber
0009|FDMS 1.0|0C|OW|1|FilmUID
0009|FDMS 1.0|F0|CS|1|BlackeningProcessFlag
0019|FDMS 1.0|90|SH|1|FilmAnnotationCharacterString1
0019|FDMS 1.0|91|SH|1|FilmAnnotationCharacterString2
0009|FDMS 1.0|05|OW|1|ImageUID
0009|FDMS 1.0|08|UL|1|ImageDisplayInformationVersionNo
0009|FDMS 1.0|09|UL|1|PatientInformationVersionNo
0009|FDMS 1.0|10|CS|1|ExposureUnitTypeCode
0009|FDMS 1.0|80|LO|1|KanjiHospitalName
0009|FDMS 1.0|90|ST|1|DistributionCode
0009|FDMS 1.0|92|SH|1|KanjiDepartmentName
0019|FDMS 1.0|15|LO|1|KanjiBodyPartForExposure
0019|FDMS 1.0|32|LO|1|KanjiMenuName
0019|FDMS 1.0|40|CS|1|ImageProcessingType
0019|FDMS 1.0|50|CS|1|EDRMode
0019|FDMS 1.0|60|SH|1|RadiographersCode
0019|FDMS 1.0|70|IS|1|SplitExposureFormat
0019|FDMS 1.0|71|IS|1|NoOfSplitExposureFrames
0019|FDMS 1.0|80|IS|1|ReadingPositionSpecification
0019|FDMS 1.0|81|IS|1|ReadingSensitivityCenter
0021|FDMS 1.0|10|CS|1|FCRImageID
0021|FDMS 1.0|30|CS|1|SetNo
0043|GEMS_PARM_01|a8|DS|3|Dual Drive Mode, Amplitude Attentuation and Phase Offset
0023|FDMS 1.0|10|SQ|1|Unknown
0023|FDMS 1.0|20|SQ|1|Unknown
0023|FDMS 1.0|30|SQ|1|Unknown
0025|FDMS 1.0|13|US|1|Unknown
0025|FDMS 1.0|15|CS|1|Unknown
0025|FDMS 1.0|20|US|2|Unknown
0025|FDMS 1.0|21|US|1|Unknown
0025|FDMS 1.0|30|US|1|Unknown
0025|FDMS 1.0|31|SS|1|Unknown
0025|FDMS 1.0|32|US|1|Unknown
0025|FDMS 1.0|33|SS|1|Unknown
0025|FDMS 1.0|34|SS|1|Unknown
0025|FDMS 1.0|40|US|1|Unknown
0025|FDMS 1.0|41|US|1|Unknown
0025|FDMS 1.0|42|US|1|Unknown
0025|FDMS 1.0|43|US|1|Unknown
0025|FDMS 1.0|50|US|1|Unknown
0025|FDMS 1.0|51|US|1|Unknown
0025|FDMS 1.0|52|US|1|Unknown
0025|FDMS 1.0|53|US|1|Unknown
0025|FDMS 1.0|60|US|1|Unknown
0025|FDMS 1.0|61|US|1|Unknown
0025|FDMS 1.0|62|US|1|Unknown
0025|FDMS 1.0|63|CS|1|Unknown
0025|FDMS 1.0|70|US|1|Unknown
0025|FDMS 1.0|71|US|1|Unknown
0025|FDMS 1.0|72|US|1|Unknown
0025|FDMS 1.0|73|US|1-n|Unknown
0025|FDMS 1.0|74|US|1-n|Unknown
0025|FDMS 1.0|80|US|1|Unknown
0025|FDMS 1.0|81|US|1|Unknown
0025|FDMS 1.0|82|US|1|Unknown
0025|FDMS 1.0|83|US|1-n|Unknown
0025|FDMS 1.0|84|US|1-n|Unknown
0025|FDMS 1.0|90|US|1|Unknown
0025|FDMS 1.0|91|US|1|Unknown
0025|FDMS 1.0|92|US|1|Unknown
0025|FDMS 1.0|93|US|1|Unknown
0025|FDMS 1.0|94|US|1|Unknown
0025|FDMS 1.0|95|US|1|Unknown
0025|FDMS 1.0|96|CS|1|Unknown
0025|FDMS 1.0|a0|US|1|Unknown
0025|FDMS 1.0|a1|SS|1|Unknown
0025|FDMS 1.0|a2|US|1|Unknown
0025|FDMS 1.0|a3|SS|1|Unknown
0027|FDMS 1.0|10|SQ|1|Unknown
0027|FDMS 1.0|20|SQ|1|Unknown
0027|FDMS 1.0|30|SQ|1|Unknown
0027|FDMS 1.0|40|SQ|1|Unknown
0027|FDMS 1.0|50|SQ|1|Unknown
0027|FDMS 1.0|60|SQ|1|Unknown
0027|FDMS 1.0|70|SQ|1|Unknown
0027|FDMS 1.0|80|SQ|1|Unknown
0027|FDMS 1.0|a0|IS|1|Unknown
0027|FDMS 1.0|a1|CS|2|Unknown
0027|FDMS 1.0|a2|CS|2|Unknown
0027|FDMS 1.0|a3|SS|1-n|Unknown
0029|FDMS 1.0|20|CS|1|ImageScanningDirection
0029|FDMS 1.0|30|CS|1|ExtendedReadingSizeValue
0029|FDMS 1.0|34|US|1|MagnificationReductionRatio
0029|FDMS 1.0|44|CS|1|LineDensityCode
0021|FDMS 1.0|50|CS|1|PairProcessingInformation
0021|FDMS 1.0|80|OB|1|EquipmentTypeSpecificInformation
0025|FDMS 1.0|10|US|1|RelativeLightEmissionAmountSk
0025|FDMS 1.0|11|US|1|TermOfCorrectionForEachIPTypeSt
0025|FDMS 1.0|12|US|1|ReadingGainGp
0029|FDMS 1.0|50|CS|1|DataCompressionCode
2011|FDMS 1.0|11|CS|1|ImagePosition SpecifyingFlag
50F1|FDMS 1.0|06|CS|1|EnergySubtractionParam
50F1|FDMS 1.0|07|CS|1|SubtractionRegistrationResult
50F1|FDMS 1.0|08|CS|1|EnergySubtractionParam2
50F1|FDMS 1.0|09|SL|1|AfinConversionCoefficient
50F1|FDMS 1.0|10|CS|1|FilmOutputFormat
50F1|FDMS 1.0|20|CS|1|ImageProcessingModificationFlag
0009|FFP DATA|01|UN|1|CRHeaderInformation
0019|GE ??? From Adantage Review CS|30|LO|1|CREDRMode
0019|GE ??? From Adantage Review CS|40|LO|1|CRLatitude
0019|GE ??? From Adantage Review CS|50|LO|1|CRGroupNumber
0019|GE ??? From Adantage Review CS|70|LO|1|CRImageSerialNumber
0019|GE ??? From Adantage Review CS|80|LO|1|CRBarCodeNumber
0019|GE ??? From Adantage Review CS|90|LO|1|CRFilmOutputExposures
0009|GEMS_ACQU_01|24|DS|1|Unknown
0009|GEMS_ACQU_01|25|US|1|Unknown
0009|GEMS_ACQU_01|3e|US|1|Unknown
0009|GEMS_ACQU_01|3f|US|1|Unknown
0009|GEMS_ACQU_01|42|US|1|Unknown
0009|GEMS_ACQU_01|43|US|1|Unknown
0009|GEMS_ACQU_01|f8|US|1|Unknown
0009|GEMS_ACQU_01|fb|IS|1|Unknown
0019|GEMS_ACQU_01|01|LT|1|Unknown
0119|MRSC|1126|ST|1|PixelMaskSource
0019|GEMS_ACQU_01|05|LT|1|Unknown
0019|GEMS_ACQU_01|06|UN|1|Unknown
0019|GEMS_ACQU_01|0e|US|1|Unknown
0019|GEMS_ACQU_01|20|DS|1|Unknown
0019|GEMS_ACQU_01|22|DS|1|Unknown
0019|GEMS_ACQU_01|2d|US|1|Unknown
0019|GEMS_ACQU_01|3a|IS|1|Unknown
0019|GEMS_ACQU_01|3b|LT|1|Unknown
0019|GEMS_ACQU_01|3c|UN|1|Unknown
0019|GEMS_ACQU_01|03|DS|1|CellNumberAtTheta
0019|GEMS_ACQU_01|04|DS|1|CellSpacing
0019|GEMS_ACQU_01|0f|DS|1|HorizontalFrameOfReference
0019|GEMS_ACQU_01|11|SS|1|SeriesContrast
0019|GEMS_ACQU_01|12|SS|1|LastPseq
0019|GEMS_ACQU_01|13|SS|1|StartNumberForBaseline
0019|GEMS_ACQU_01|14|SS|1|End NumberForBaseline
0019|GEMS_ACQU_01|15|SS|1|StartNumberForEnhancedScans
0019|GEMS_ACQU_01|16|SS|1|EndNumberForEnhancedScans
0019|GEMS_ACQU_01|17|SS|1|SeriesPlane
0019|GEMS_ACQU_01|18|LO|1|FirstScanRAS
0019|GEMS_ACQU_01|19|DS|1|FirstScanLocation
0019|GEMS_ACQU_01|1a|LO|1|LastScanRAS
0019|GEMS_ACQU_01|1b|DS|1|LastScanLocation
0019|GEMS_ACQU_01|1e|DS|1|DisplayFieldOfView
0019|GEMS_ACQU_01|23|DS|1|TableSpeed
0019|GEMS_ACQU_01|24|DS|1|MidScanTime
0019|GEMS_ACQU_01|26|SL|1|DegreesOfAzimuth
0019|GEMS_ACQU_01|27|DS|1|GantryPeriod
0019|GEMS_ACQU_01|2a|DS|1|XrayOnPosition
0019|GEMS_ACQU_01|2b|DS|1|XrayOffPosition
0019|GEMS_ACQU_01|2c|SL|1|NumberOfTriggers
0019|GEMS_ACQU_01|2e|DS|1|AngleOfFirstView
0019|GEMS_ACQU_01|2f|DS|1|TriggerFrequency
0019|GEMS_ACQU_01|39|SS|1|ScanFOVType
0019|GEMS_ACQU_01|3e|UN|1|Unknown
0019|GEMS_ACQU_01|3f|UN|1|Unknown
0119|MRSC|1130|DS|1-n|UpperFitLimit
0019|GEMS_ACQU_01|48|US|1|Unknown
0019|GEMS_ACQU_01|49|US|1|Unknown
0019|GEMS_ACQU_01|54|UN|1|Unknown
0019|GEMS_ACQU_01|5d|US|1|Unknown
0019|GEMS_ACQU_01|82|US|1|Unknown
0019|GEMS_ACQU_01|83|DS|1|Unknown
0019|GEMS_ACQU_01|86|US|1|Unknown
0019|GEMS_ACQU_01|99|US|1|Unknown
0019|GEMS_ACQU_01|42|SS|1|SegmentNumber
0019|GEMS_ACQU_01|43|SS|1|TotalSegmentsRequested
0019|GEMS_ACQU_01|44|DS|1|InterscanDelay
0019|GEMS_ACQU_01|47|SS|1|ViewCompressionFactor
0019|GEMS_ACQU_01|4a|SS|1|TotalNumberOfRefChannels
0019|GEMS_ACQU_01|4b|SL|1|DataSizeForScanData
0019|GEMS_ACQU_01|52|SS|1|ReconPostProcessingFlag
0019|GEMS_ACQU_01|57|SS|1|CTWaterNumber
0019|GEMS_ACQU_01|58|SS|1|CTBoneNumber
0019|GEMS_ACQU_01|5a|FL|1|AcquisitionDuration
0019|GEMS_ACQU_01|5e|SL|1|NumberOfChannels1To512
0019|GEMS_ACQU_01|5f|SL|1|IncrementBetweenChannels
0019|GEMS_ACQU_01|60|SL|1|StartingView
0019|GEMS_ACQU_01|61|SL|1|NumberOfViews
0019|GEMS_ACQU_01|62|SL|1|IncrementBetweenViews
0019|GEMS_ACQU_01|6b|SS|1|FieldOfViewInDetectorCells
0019|GEMS_ACQU_01|70|SS|1|ValueOfBackProjectionButton
0019|GEMS_ACQU_01|71|SS|1|SetIfFatqEstimatesWereUsed
0019|GEMS_ACQU_01|72|DS|1|ZChannelAvgOverViews
0019|GEMS_ACQU_01|73|DS|1|AvgOfLeftRefChannelsOverViews
0019|GEMS_ACQU_01|74|DS|1|MaxLeftChannelOverViews
0019|GEMS_ACQU_01|75|DS|1|AvgOfRightRefChannelsOverViews
0019|GEMS_ACQU_01|76|DS|1|MaxRightChannelOverViews
0019|GEMS_ACQU_01|7d|DS|1|SecondEcho
0019|GEMS_ACQU_01|7e|SS|1|NumberOfEchos
0019|GEMS_ACQU_01|7f|DS|1|TableDelta
0019|GEMS_ACQU_01|81|SS|1|Contiguous
0019|GEMS_ACQU_01|84|DS|1|PeakSAR
0019|GEMS_ACQU_01|85|SS|1|MonitorSAR
0019|GEMS_ACQU_01|87|DS|1|CardiacRepetition Time
0019|GEMS_ACQU_01|88|SS|1|ImagesPerCardiacCycle
0019|GEMS_ACQU_01|8a|SS|1|ActualReceiveGainAnalog
0019|GEMS_ACQU_01|8b|SS|1|ActualReceiveGainDigital
0019|GEMS_ACQU_01|8d|DS|1|DelayAfterTrigger
0019|GEMS_ACQU_01|8f|SS|1|SwapPhaseFrequency
0019|GEMS_ACQU_01|90|SS|1|PauseInterval
0019|GEMS_ACQU_01|91|DS|1|PulseTime
0019|GEMS_ACQU_01|93|DS|1|CenterFrequency
0019|GEMS_ACQU_01|94|SS|1|TransmitGain
0019|GEMS_ACQU_01|95|SS|1|AnalogReceiverGain
0019|GEMS_ACQU_01|96|SS|1|DigitalReceiverGain
0019|GEMS_ACQU_01|97|SL|1|BitmapDefiningCVs
0019|GEMS_ACQU_01|98|SS|1|CenterFrequencyMethod
0019|GEMS_ACQU_01|9b|SS|1|PulseSequenceMode
0019|GEMS_ACQU_01|9c|LO|1|PulseSequenceName
0019|GEMS_ACQU_01|9d|DT|1|PulseSequenceDate
0019|GEMS_ACQU_01|d4|US|1|Unknown
0019|GEMS_ACQU_01|9f|SS|1|TransmittingCoil
0019|GEMS_ACQU_01|a0|SS|1|SurfaceCoilType
0019|GEMS_ACQU_01|a1|SS|1|ExtremityCoilFlag
0019|GEMS_ACQU_01|a2|SL|1|RawDataRunNumber
0019|GEMS_ACQU_01|a3|UL|1|CalibratedFieldStrength
0019|GEMS_ACQU_01|a4|SS|1|SATFatWaterBone
0019|GEMS_ACQU_01|a5|DS|1|ReceiveBandwidth
0019|GEMS_ACQU_01|a7|DS|1|UserData
0019|GEMS_ACQU_01|a8|DS|1|UserData
0019|GEMS_ACQU_01|a9|DS|1|UserData
0019|GEMS_ACQU_01|aa|DS|1|UserData
0019|GEMS_ACQU_01|ab|DS|1|UserData
0019|GEMS_ACQU_01|ac|DS|1|UserData
0019|GEMS_ACQU_01|ad|DS|1|UserData
0019|GEMS_ACQU_01|ae|DS|1|UserData
0019|GEMS_ACQU_01|af|DS|1|UserData
0019|GEMS_ACQU_01|b0|DS|1|UserData
0019|GEMS_ACQU_01|b1|DS|1|UserData
0019|GEMS_ACQU_01|b3|DS|1|UserData
0019|GEMS_ACQU_01|b4|DS|1|UserData
0019|GEMS_ACQU_01|b5|DS|1|UserData
0019|GEMS_ACQU_01|b6|DS|1|UserData
0019|GEMS_ACQU_01|b7|DS|1|UserData
0019|GEMS_ACQU_01|b8|DS|1|UserData
0019|GEMS_ACQU_01|b9|DS|1|UserData
0019|GEMS_ACQU_01|ba|DS|1|UserData
0019|GEMS_ACQU_01|bb|DS|1|UserData
0019|GEMS_ACQU_01|bc|DS|1|UserData
0019|GEMS_ACQU_01|bd|DS|1|UserData
0019|GEMS_ACQU_01|be|DS|1|ProjectionAngle
0019|GEMS_ACQU_01|c0|SS|1|SaturationPlanes
0019|GEMS_ACQU_01|c1|SS|1|SurfaceCoilIntensityCorrectionFlag
0019|GEMS_ACQU_01|c2|SS|1|SATLocationR
0019|GEMS_ACQU_01|c3|SS|1|SATLocationL
0019|GEMS_ACQU_01|c4|SS|1|SATLocationA
0019|GEMS_ACQU_01|c5|SS|1|SATLocationP
0019|GEMS_ACQU_01|c6|SS|1|SATLocationH
0019|GEMS_ACQU_01|c7|SS|1|SATLocationF
0019|GEMS_ACQU_01|c8|SS|1|SATThicknessRL
0019|GEMS_ACQU_01|c9|SS|1|SATThicknessAP
0019|GEMS_ACQU_01|ca|SS|1|SATThicknessHF
0019|GEMS_ACQU_01|cc|SS|1|VelocityEncoding
0019|GEMS_ACQU_01|cd|SS|1|ThicknessDisclaimer
0019|GEMS_ACQU_01|ce|SS|1|PrescanType
0019|GEMS_ACQU_01|cf|SS|1|PrescanStatus
0019|GEMS_ACQU_01|d0|SH|1|RawDataType
0019|GEMS_ACQU_01|d2|SS|1|ProjectionAlgorithm
0019|GEMS_ACQU_01|d3|SH|1|ProjectionAlgorithm
0019|GEMS_ACQU_01|d5|SS|1|FractionalEcho
0019|GEMS_ACQU_01|d6|SS|1|PrepPulse
0019|GEMS_ACQU_01|d7|SS|1|CardiacPhases
0019|GEMS_ACQU_01|d8|SS|1|VariableEchoFlag
0019|GEMS_ACQU_01|d9|DS|1|ConcatenatedSAT
0019|GEMS_ACQU_01|da|SS|1|ReferenceChannelUsed
0019|GEMS_ACQU_01|db|DS|1|BackProjectorCoefficient
0019|GEMS_ACQU_01|dc|SS|1|PrimarySpeedCorrectionUsed
0119|MRSC|1131|DS|1-n|LowerFitLimit
0019|GEMS_ACQU_01|e1|DS|1|Unknown
0019|GEMS_ACQU_01|e3|LT|1|Unknown
0019|GEMS_ACQU_01|e4|LT|1|Unknown
0019|GEMS_ACQU_01|e5|IS|1|Unknown
0019|GEMS_ACQU_01|e6|US|1|Unknown
0019|GEMS_ACQU_01|e8|DS|1|Unknown
0019|GEMS_ACQU_01|e9|DS|1|Unknown
0019|GEMS_ACQU_01|eb|DS|1|Unknown
0019|GEMS_ACQU_01|ec|US|1|Unknown
0019|GEMS_ACQU_01|f0|UN|1|Unknown
0019|GEMS_ACQU_01|f1|LT|1|Unknown
0019|GEMS_ACQU_01|f3|LT|1|Unknown
0019|GEMS_ACQU_01|f4|LT|1|Unknown
0023|GEMS_ACRQA_1.0 BLOCK1|00|LO|1|CRExposureMenuCode
0023|GEMS_ACRQA_1.0 BLOCK1|10|LO|1|CRExposureMenuString
0023|GEMS_ACRQA_1.0 BLOCK1|20|LO|1|CREDRMode
0023|GEMS_ACRQA_1.0 BLOCK1|30|LO|1|CRLatitude
0023|GEMS_ACRQA_1.0 BLOCK1|40|LO|1|CRGroupNumber
0023|GEMS_ACRQA_1.0 BLOCK1|50|US|1|CRImageSerialNumber
0023|GEMS_ACRQA_1.0 BLOCK1|60|LO|1|CRBarCodeNumber
0023|GEMS_ACRQA_1.0 BLOCK1|70|LO|1|CRFilmOutputExposure
0023|GEMS_ACRQA_1.0 BLOCK1|80|LO|1|CRFilmFormat
0023|GEMS_ACRQA_1.0 BLOCK1|90|LO|1|CRSShiftString
0023|GEMS_ACRQA_1.0 BLOCK2|00|US|1|CRSShift
0023|GEMS_ACRQA_1.0 BLOCK2|10|DS|1|CRCShift
0023|GEMS_ACRQA_1.0 BLOCK2|20|DS|1|CRGT
0023|GEMS_ACRQA_1.0 BLOCK2|30|DS|1|CRGA
0023|GEMS_ACRQA_1.0 BLOCK2|40|DS|1|CRGC
0023|GEMS_ACRQA_1.0 BLOCK2|50|DS|1|CRGS
0023|GEMS_ACRQA_1.0 BLOCK2|60|DS|1|CRRT
0023|GEMS_ACRQA_1.0 BLOCK2|70|DS|1|CRRE
0023|GEMS_ACRQA_1.0 BLOCK2|80|US|1|CRRN
0023|GEMS_ACRQA_1.0 BLOCK2|90|DS|1|CRDRT
0023|GEMS_ACRQA_1.0 BLOCK3|00|DS|1|CRDRE
0023|GEMS_ACRQA_1.0 BLOCK3|10|US|1|CRDRN
0023|GEMS_ACRQA_1.0 BLOCK3|20|DS|1|CRORE
0023|GEMS_ACRQA_1.0 BLOCK3|30|US|1|CRORN
0023|GEMS_ACRQA_1.0 BLOCK3|40|US|1|CRORD
0023|GEMS_ACRQA_1.0 BLOCK3|50|LO|1|CRCassetteSize
0023|GEMS_ACRQA_1.0 BLOCK3|60|LO|1|CRMachineID
0023|GEMS_ACRQA_1.0 BLOCK3|70|LO|1|CRMachineType
0023|GEMS_ACRQA_1.0 BLOCK3|80|LO|1|CRTechnicianCode
0023|GEMS_ACRQA_1.0 BLOCK3|90|LO|1|CREnergySubtractionParameters
0023|GEMS_ACRQA_2.0 BLOCK1|00|LO|1|CRExposureMenuCode
0023|GEMS_ACRQA_2.0 BLOCK1|10|LO|1|CRExposureMenuString
0023|GEMS_ACRQA_2.0 BLOCK1|20|LO|1|CREDRMode
0023|GEMS_ACRQA_2.0 BLOCK1|30|LO|1|CRLatitude
0023|GEMS_ACRQA_2.0 BLOCK1|40|LO|1|CRGroupNumber
0019|GEMS_ACQU_01|de|DS|1|DynamicZAlphaValue
0019|GEMS_ACQU_01|df|DS|1|UserData
0019|GEMS_ACQU_01|e0|DS|1|UserData
0019|GEMS_ACQU_01|e2|DS|1|VelocityEncodeScale
0019|GEMS_ACQU_01|f2|SS|1|FastPhases
0019|GEMS_ACQU_01|f9|DS|1|TransmissionGain
0023|GEMS_ACRQA_2.0 BLOCK1|50|US|1|CRImageSerialNumber
0023|GEMS_ACRQA_2.0 BLOCK1|60|LO|1|CRBarCodeNumber
0023|GEMS_ACRQA_2.0 BLOCK1|70|LO|1|CRFilmOutputExposure
0023|GEMS_ACRQA_2.0 BLOCK1|80|LO|1|CRFilmFormat
0023|GEMS_ACRQA_2.0 BLOCK1|90|LO|1|CRSShiftString
0023|GEMS_ACRQA_2.0 BLOCK2|00|US|1|CRSShift
0023|GEMS_ACRQA_2.0 BLOCK2|10|LO|1|CRCShift
0023|GEMS_ACRQA_2.0 BLOCK2|20|LO|1|CRGT
0023|GEMS_ACRQA_2.0 BLOCK2|30|DS|1|CRGA
0023|GEMS_ACRQA_2.0 BLOCK2|40|DS|1|CRGC
0023|GEMS_ACRQA_2.0 BLOCK2|50|DS|1|CRGS
0023|GEMS_ACRQA_2.0 BLOCK2|60|LO|1|CRRT
0023|GEMS_ACRQA_2.0 BLOCK2|70|DS|1|CRRE
0023|GEMS_ACRQA_2.0 BLOCK2|80|US|1|CRRN
0023|GEMS_ACRQA_2.0 BLOCK2|90|DS|1|CRDRT
0023|GEMS_ACRQA_2.0 BLOCK3|00|DS|1|CRDRE
0023|GEMS_ACRQA_2.0 BLOCK3|10|US|1|CRDRN
0023|GEMS_ACRQA_2.0 BLOCK3|20|DS|1|CRORE
0023|GEMS_ACRQA_2.0 BLOCK3|30|US|1|CRORN
0023|GEMS_ACRQA_2.0 BLOCK3|40|US|1|CRORD
0023|GEMS_ACRQA_2.0 BLOCK3|50|LO|1|CRCassetteSize
0023|GEMS_ACRQA_2.0 BLOCK3|60|LO|1|CRMachineID
0023|GEMS_ACRQA_2.0 BLOCK3|70|LO|1|CRMachineType
0023|GEMS_ACRQA_2.0 BLOCK3|80|LO|1|CRTechnicianCode
0023|GEMS_ACRQA_2.0 BLOCK3|90|LO|1|CREnergySubtractionParameters
0023|GEMS_ACRQA_2.0 BLOCK3|f0|LO|1|CRDistributionCode
0023|GEMS_ACRQA_2.0 BLOCK3|ff|US|1|CRShuttersApplied
0047|GEMS_ADWSoft_3D1|01|SQ|1|Reconstruction Parameters Sequence
0047|GEMS_ADWSoft_3D1|50|UL|1|VolumeVoxelCount
0047|GEMS_ADWSoft_3D1|51|UL|1|VolumeSegmentCount
0047|GEMS_ADWSoft_3D1|53|US|1|VolumeSliceSize
0047|GEMS_ADWSoft_3D1|54|US|1|VolumeSliceCount
0047|GEMS_ADWSoft_3D1|55|SL|1|VolumeThresholdValue
0047|GEMS_ADWSoft_3D1|57|DS|1|VolumeVoxelRatio
0047|GEMS_ADWSoft_3D1|58|DS|1|VolumeVoxelSize
0047|GEMS_ADWSoft_3D1|59|US|1|VolumeZPositionSize
0047|GEMS_ADWSoft_3D1|60|DS|9|VolumeBaseLine
0047|GEMS_ADWSoft_3D1|61|DS|3|VolumeCenterPoint
0047|GEMS_ADWSoft_3D1|63|SL|1|VolumeSkewBase
0047|GEMS_ADWSoft_3D1|64|DS|9|VolumeRegistrationTransformRotationMatrix
0047|GEMS_ADWSoft_3D1|65|DS|3|VolumeRegistrationTransformTranslationVector
0047|GEMS_ADWSoft_3D1|70|DS|1-n|KVPList
0047|GEMS_ADWSoft_3D1|71|IS|1-n|XRayTubeCurrentList
0047|GEMS_ADWSoft_3D1|72|IS|1-n|ExposureList
0047|GEMS_ADWSoft_3D1|80|LO|1|AcquisitionDLXIdentifier
0047|GEMS_ADWSoft_3D1|85|SQ|1|AcquisitionDLX2DSeriesSequence
0047|GEMS_ADWSoft_3D1|89|DS|1-n|ContrastAgentVolumeList
0047|GEMS_ADWSoft_3D1|8A|US|1|NumberOfInjections
0047|GEMS_ADWSoft_3D1|8B|US|1|FrameCount
0047|GEMS_ADWSoft_3D1|91|LO|1|XA3DReconstructionAlgorithmName
0047|GEMS_ADWSoft_3D1|92|CS|1|XA3DReconstructionAlgorithmVersion
0047|GEMS_ADWSoft_3D1|93|DA|1|DLXCalibrationDate
0047|GEMS_ADWSoft_3D1|94|TM|1|DLXCalibrationTime
0047|GEMS_ADWSoft_3D1|95|CS|1|DLXCalibrationStatus
0047|GEMS_ADWSoft_3D1|96|IS|1-n|UsedFrames
0047|GEMS_ADWSoft_3D1|98|US|1|TransformCount
0047|GEMS_ADWSoft_3D1|99|SQ|1|TransformSequence
0047|GEMS_ADWSoft_3D1|9A|DS|9|TransformRotationMatrix
0047|GEMS_ADWSoft_3D1|9B|DS|3|TransformTranslationVector
0047|GEMS_ADWSoft_3D1|9C|LO|1|TransformLabel
0047|GEMS_ADWSoft_3D1|B0|SQ|1|WireframeList
0047|GEMS_ADWSoft_3D1|B1|US|1|WireframeCount
0047|GEMS_ADWSoft_3D1|B2|US|1|LocationSystem
0047|GEMS_ADWSoft_3D1|B5|LO|1|WireframeName
0047|GEMS_ADWSoft_3D1|B6|LO|1|WireframeGroupName
0047|GEMS_ADWSoft_3D1|B7|LO|1|WireframeColor
0047|GEMS_ADWSoft_3D1|B8|SL|1|WireframeAttributes
0047|GEMS_ADWSoft_3D1|B9|SL|1|WireframePointCount
0047|GEMS_ADWSoft_3D1|BA|SL|1|WireframeTimestamp
0047|GEMS_ADWSoft_3D1|BB|SQ|1|WireframePointList
0047|GEMS_ADWSoft_3D1|BC|DS|3|WireframePointsCoordinates
0047|GEMS_ADWSoft_3D1|C0|DS|3|VolumeUpperLeftHighCornerRAS
0047|GEMS_ADWSoft_3D1|C1|DS|9|VolumeSliceToRASRotationMatrix
0047|GEMS_ADWSoft_3D1|C2|DS|1|VolumeUpperLeftHighCornerTLOC
0047|GEMS_ADWSoft_3D1|D1|OB|1|VolumeSegmentList
0047|GEMS_ADWSoft_3D1|D2|OB|1|VolumeGradientList
0047|GEMS_ADWSoft_3D1|D3|OB|1|VolumeDensityList
0047|GEMS_ADWSoft_3D1|D4|OB|1|VolumeZPositionList
0047|GEMS_ADWSoft_3D1|D5|OB|1|VolumeOriginalIndexList
0039|GEMS_ADWSoft_DPO|80|IS|1|PrivateEntityNumber
0039|GEMS_ADWSoft_DPO|85|DA|1|PrivateEntityDate
0039|GEMS_ADWSoft_DPO|90|TM|1|PrivateEntityTime
0039|GEMS_ADWSoft_DPO|95|LO|1|PrivateEntityLaunchCommand
0039|GEMS_ADWSoft_DPO|AA|CS|1|PrivateEntityType
0033|GEMS_CTHD_01|02|UN|1|Unknown
0037|GEMS_DRS_1|10|LO|1|ReferringDepartment
0037|GEMS_DRS_1|20|US|1|ScreenNumber
0037|GEMS_DRS_1|40|SH|1|LeftOrientation
0037|GEMS_DRS_1|42|SH|1|RightOrientation
0037|GEMS_DRS_1|50|CS|1|Inversion
0037|GEMS_DRS_1|60|US|1|DSA
0009|GEMS_GENIE_1|10|LO|1|Unknown
0009|GEMS_GENIE_1|11|SL|1|StudyFlags
0009|GEMS_GENIE_1|12|SL|1|StudyType
0009|GEMS_GENIE_1|1e|UI|1|Unknown
0009|GEMS_GENIE_1|20|LO|1|Unknown
0009|GEMS_GENIE_1|21|SL|1|SeriesFlags
0009|GEMS_GENIE_1|22|SH|1|UserOrientation
0009|GEMS_GENIE_1|23|SL|1|InitiationType
0009|GEMS_GENIE_1|24|SL|1|InitiationDelay
0009|GEMS_GENIE_1|25|SL|1|InitiationCountRate
0009|GEMS_GENIE_1|26|SL|1|NumberEnergySets
0009|GEMS_GENIE_1|27|SL|1|NumberDetectors
0009|GEMS_GENIE_1|29|SL|1|Unknown
0009|GEMS_GENIE_1|2a|SL|1|Unknown
0009|GEMS_GENIE_1|2c|LO|1|SeriesComments
0009|GEMS_GENIE_1|2d|SL|1|TrackBeatAverage
0009|GEMS_GENIE_1|2e|FD|1|DistancePrescribed
0009|GEMS_GENIE_1|30|LO|1|Unknown
0009|GEMS_GENIE_1|35|SL|1|GantryLocusType
0009|GEMS_GENIE_1|37|SL|1|StartingHeartRate
0009|GEMS_GENIE_1|38|SL|1|RRWindowWidth
0009|GEMS_GENIE_1|39|SL|1|RRWindowOffset
0009|GEMS_GENIE_1|3a|SL|1|PercentCycleImaged
0009|GEMS_GENIE_1|40|LO|1|Unknown
0009|GEMS_GENIE_1|41|SL|1|PatientFlags
0009|GEMS_GENIE_1|42|DA|1|PatientCreationDate
0009|GEMS_GENIE_1|43|TM|1|PatientCreationTime
0011|GEMS_GENIE_1|0a|SL|1|SeriesType
0011|GEMS_GENIE_1|0b|SL|1|EffectiveSeriesDuration
0011|GEMS_GENIE_1|0c|SL|1|NumBeats
0011|GEMS_GENIE_1|0d|LO|1|RadioNuclideName
0011|GEMS_GENIE_1|10|LO|1|Unknown
0011|GEMS_GENIE_1|12|LO|1|DatasetName
0011|GEMS_GENIE_1|13|SL|1|DatasetType
0011|GEMS_GENIE_1|15|SL|1|DetectorNumber
0011|GEMS_GENIE_1|16|SL|1|EnergyNumber
0011|GEMS_GENIE_1|17|SL|1|RRIntervalWindowNumber
0011|GEMS_GENIE_1|18|SL|1|MGBinNumber
0011|GEMS_GENIE_1|19|FD|1|RadiusOfRotation
0011|GEMS_GENIE_1|1a|SL|1|DetectorCountZone
0011|GEMS_GENIE_1|1b|SL|1|NumEnergyWindows
0011|GEMS_GENIE_1|1c|SL|4|EnergyOffset
0011|GEMS_GENIE_1|1d|SL|1|EnergyRange
0011|GEMS_GENIE_1|1f|SL|1|ImageOrientation
0011|GEMS_GENIE_1|23|SL|1|UseFOVMask
0011|GEMS_GENIE_1|24|SL|1|FOVMaskYCutoffAngle
0011|GEMS_GENIE_1|25|SL|1|FOVMaskCutoffAngle
0011|GEMS_GENIE_1|26|SL|1|TableOrientation
0011|GEMS_GENIE_1|27|SL|2|ROITopLeft
0011|GEMS_GENIE_1|28|SL|2|ROIBottomRight
0011|GEMS_GENIE_1|30|LO|1|Unknown
0011|GEMS_GENIE_1|33|LO|1|EnergyCorrectName
0011|GEMS_GENIE_1|34|LO|1|SpatialCorrectName
0011|GEMS_GENIE_1|35|LO|1|TuningCalibName
0011|GEMS_GENIE_1|36|LO|1|UniformityCorrectName
0011|GEMS_GENIE_1|37|LO|1|AcquisitionSpecificCorrectName
0011|GEMS_GENIE_1|38|SL|1|ByteOrder
0011|GEMS_GENIE_1|3a|SL|1|PictureFormat
0011|GEMS_GENIE_1|3b|FD|1|PixelScale
0011|GEMS_GENIE_1|3c|FD|1|PixelOffset
0011|GEMS_GENIE_1|3e|SL|1|FOVShape
0011|GEMS_GENIE_1|3f|SL|1|DatasetFlags
0011|GEMS_GENIE_1|44|FD|1|ThresholdCenter
0011|GEMS_GENIE_1|45|FD|1|ThresholdWidth
0011|GEMS_GENIE_1|46|SL|1|InterpolationType
0011|GEMS_GENIE_1|55|FD|1|Period
0011|GEMS_GENIE_1|56|FD|1|ElapsedTime
0013|GEMS_GENIE_1|10|FD|2|DigitalFOV
0013|GEMS_GENIE_1|11|SL|1|Unknown
0013|GEMS_GENIE_1|12|SL|1|Unknown
0013|GEMS_GENIE_1|16|SL|1|AutoTrackPeak
0013|GEMS_GENIE_1|17|SL|1|AutoTrackWidth
0013|GEMS_GENIE_1|18|FD|1|TransmissionScanTime
0013|GEMS_GENIE_1|19|FD|1|TransmissionMaskWidth
0013|GEMS_GENIE_1|1a|FD|1|CopperAttenuatorThickness
0013|GEMS_GENIE_1|1c|FD|1|Unknown
0013|GEMS_GENIE_1|1d|FD|1|Unknown
0013|GEMS_GENIE_1|1e|FD|1-n|TomoViewOffset
0013|GEMS_GENIE_1|26|LT|1|StudyComments
0033|GEMS_GNHD_01|01|UN|1|Unknown
0033|GEMS_GNHD_01|02|UN|1|Unknown
0119|MRSC|1140|LO|1|GradientMatrixMethod
0009|GEMS_IDEN_01|e8|UL|1|Unknown
0009|GEMS_IDEN_01|02|SH|1|SuiteId
0009|GEMS_IDEN_01|04|SH|1|ProductId
0009|GEMS_IDEN_01|17|LT|1|Unknown
0009|GEMS_IDEN_01|1a|US|1|Unknown
0009|GEMS_IDEN_01|20|US|1|Unknown
0009|GEMS_IDEN_01|27|SL|1|ImageActualDate
0009|GEMS_IDEN_01|2f|LT|1|Unknown
0009|GEMS_IDEN_01|30|SH|1|ServiceId
0009|GEMS_IDEN_01|31|SH|1|MobileLocationNumber
0009|GEMS_IDEN_01|e2|LT|1|Unknown
0009|GEMS_IDEN_01|e3|UI|1|EquipmentUID
0009|GEMS_IDEN_01|e6|SH|1|GenesisVersionNow
0009|GEMS_IDEN_01|e7|UL|1|ExamRecordChecksum
0009|GEMS_IDEN_01|e9|SL|1|ActualSeriesDataTimeStamp
0027|GEMS_IMAG_01|06|SL|1|ImageArchiveFlag
0027|GEMS_IMAG_01|10|SS|1|ScoutType
0027|GEMS_IMAG_01|1d|SS|1|VmaPhase
0027|GEMS_IMAG_01|1e|SL|1|VmaMod
0027|GEMS_IMAG_01|1f|SL|1|VmaClip
0027|GEMS_IMAG_01|20|SS|1|SmartScanOnOffFlag
0027|GEMS_IMAG_01|30|SH|1|ForeignImageRevision
0027|GEMS_IMAG_01|31|SS|1|ImagingMode
0027|GEMS_IMAG_01|32|SS|1|PulseSequence
0027|GEMS_IMAG_01|33|SL|1|ImagingOptions
0027|GEMS_IMAG_01|35|SS|1|PlaneType
0027|GEMS_IMAG_01|36|SL|1|ObliquePlane
0027|GEMS_IMAG_01|40|SH|1|RASLetterOfImageLocation
0027|GEMS_IMAG_01|41|FL|1|ImageLocation
0027|GEMS_IMAG_01|42|FL|1|CenterRCoordOfPlaneImage
0027|GEMS_IMAG_01|43|FL|1|CenterACoordOfPlaneImage
0027|GEMS_IMAG_01|45|FL|1|NormalRCoord
0027|GEMS_IMAG_01|46|FL|1|NormalACoord
0027|GEMS_IMAG_01|47|FL|1|NormalSCoord
0027|GEMS_IMAG_01|48|FL|1|RCoordOfTopRightCorner
0027|GEMS_IMAG_01|49|FL|1|ACoordOfTopRightCorner
0027|GEMS_IMAG_01|4a|FL|1|SCoordOfTopRightCorner
0027|GEMS_IMAG_01|4b|FL|1|RCoordOfBottomRightCorner
0027|GEMS_IMAG_01|4c|FL|1|ACoordOfBottomRightCorner
0027|GEMS_IMAG_01|4d|FL|1|SCoordOfBottomRightCorner
0027|GEMS_IMAG_01|50|FL|1|TableStartLocation
0027|GEMS_IMAG_01|51|FL|1|TableEndLocation
0027|GEMS_IMAG_01|52|SH|1|RASLetterForSideOfImage
0027|GEMS_IMAG_01|53|SH|1|RASLetterForAnteriorPosterior
0027|GEMS_IMAG_01|54|SH|1|RASLetterForScoutStartLoc
0027|GEMS_IMAG_01|55|SH|1|RASLetterForScoutEndLoc
0027|GEMS_IMAG_01|60|FL|1|ImageDimensionX
0027|GEMS_IMAG_01|61|FL|1|ImageDimensionY
0027|GEMS_IMAG_01|62|FL|1|NumberOfExcitations
0029|GEMS_IMPS_01|04|SL|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|05|DS|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|07|SL|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|08|SH|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|09|SH|1|LowerRangeOfPixels
0119|MRSC|1141|DS|1-n|GradientMatrix
0029|GEMS_IMPS_01|15|SL|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|16|SL|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|17|SL|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|18|SL|1|UpperRangeOfPixels
0029|GEMS_IMPS_01|1a|SL|1|LengthOfTotalHeaderInBytes
0029|GEMS_IMPS_01|26|SS|1|VersionOfHeaderStructure
0029|GEMS_IMPS_01|34|SL|1|AdvantageCompOverflow
0029|GEMS_IMPS_01|35|SL|1|AdvantageCompUnderflow
0043|GEMS_PARM_01|01|SS|1|BitmapOfPrescanOptions
0043|GEMS_PARM_01|02|SS|1|GradientOffsetInX
0043|GEMS_PARM_01|04|SS|1|GradientOffsetInZ
0043|GEMS_PARM_01|05|SS|1|ImageIsOriginalOrUnoriginal
0043|GEMS_PARM_01|06|SS|1|NumberOfEPIShots
0043|GEMS_PARM_01|07|SS|1|ViewsPerSegment
0043|GEMS_PARM_01|08|SS|1|RespiratoryRateInBPM
0043|GEMS_PARM_01|09|SS|1|RespiratoryTriggerPoint
0043|GEMS_PARM_01|0a|SS|1|TypeOfReceiverUsed
0043|GEMS_PARM_01|0b|DS|1|PeakRateOfChangeOfGradientField
0043|GEMS_PARM_01|0c|DS|1|LimitsInUnitsOfPercent
0043|GEMS_PARM_01|0d|DS|1|PSDEstimatedLimit
0043|GEMS_PARM_01|0e|DS|1|PSDEstimatedLimitInTeslaPerSecond
0043|GEMS_PARM_01|0f|DS|1|SARAvgHead
0043|GEMS_PARM_01|10|US|1|WindowValue
0043|GEMS_PARM_01|11|US|1|TotalInputViews
0043|GEMS_PARM_01|12|SS|3|XrayChain
0043|GEMS_PARM_01|13|SS|5|ReconKernelParameters
0043|GEMS_PARM_01|14|SS|3|CalibrationParameters
0043|GEMS_PARM_01|15|SS|3|TotalOutputViews
0043|GEMS_PARM_01|16|SS|5|NumberOfOverranges
0043|GEMS_PARM_01|18|DS|3|BBH Coefficients
0043|GEMS_PARM_01|19|SS|1|NumberOfBBHChainsToBlend
0043|GEMS_PARM_01|1a|SL|1|StartingChannelNumber
0043|GEMS_PARM_01|1b|SS|1|PPScanParameters
0043|GEMS_PARM_01|1c|SS|1|GEImageIntegrity
0043|GEMS_PARM_01|1d|SS|1|LevelValue
0043|GEMS_PARM_01|1e|DS|1|DeltaStartTime
0043|GEMS_PARM_01|1f|SL|1|MaxOverrangesInAView
0043|GEMS_PARM_01|20|DS|1|AvgOverrangesAllViews
0043|GEMS_PARM_01|21|SS|1|CorrectedAfterglowTerms
0043|GEMS_PARM_01|25|SS|6|ReferenceChannels
0043|GEMS_PARM_01|26|US|6|NoViewsRefChannelsBlocked
0043|GEMS_PARM_01|27|SH|1|ScanPitchRatio
0043|GEMS_PARM_01|28|OB|1|UniqueImageIdentifier
0043|GEMS_PARM_01|29|OB|1|HistogramTables
0043|GEMS_PARM_01|2a|OB|1|UserDefinedData
0043|GEMS_PARM_01|2b|SS|4|PrivateScanOptions
0043|GEMS_PARM_01|2c|SS|1|EffectiveEchoSpacing
0043|GEMS_PARM_01|2e|SH|1|StringSlopField2
0043|GEMS_PARM_01|2f|SS|1|RawDataType
0043|GEMS_PARM_01|30|SS|1|RawDataType
0043|GEMS_PARM_01|31|DS|2|RACoordOfTargetReconCentre
0043|GEMS_PARM_01|32|SS|1|RawDataType
0043|GEMS_PARM_01|33|FL|1|NegScanSpacing
0043|GEMS_PARM_01|34|IS|1|OffsetFrequency
0043|GEMS_PARM_01|35|UL|1|UserUsageTag
0119|MRSC|1180|SQ|1|FitMapSQ
0021|GEMS_RELA_01|15|US|1|Unknown
0021|GEMS_RELA_01|16|SS|1|Unknown
0021|GEMS_RELA_01|4e|US|1|Unknown
0021|GEMS_RELA_01|70|LT|1|Unknown
0021|GEMS_RELA_01|71|LT|1|Unknown
0019|SIEMENS RA GEN|52|SS|1|TableTilt
0021|GEMS_RELA_01|05|SH|1|GenesisVersionNow
0021|GEMS_RELA_01|07|UL|1|SeriesRecordChecksum
0021|GEMS_RELA_01|18|SH|1|GenesisVersionNow
0021|GEMS_RELA_01|19|UL|1|AcqReconRecordChecksum
0021|GEMS_RELA_01|20|DS|1|TableStartLocation
0021|GEMS_RELA_01|35|SS|1|SeriesFromWhichPrescribed
0021|GEMS_RELA_01|36|SS|1|ImageFromWhichPrescribed
0021|GEMS_RELA_01|37|SS|1|ScreenFormat
0021|GEMS_RELA_01|4a|LO|1|AnatomicalReferenceForScout
0021|GEMS_RELA_01|4f|SS|1|LocationsInAcquisition
0021|GEMS_RELA_01|50|SS|1|GraphicallyPrescribed
0021|GEMS_RELA_01|51|DS|1|RotationFromSourceXRot
0021|GEMS_RELA_01|52|DS|1|RotationFromSourceYRot
0021|GEMS_RELA_01|53|DS|1|RotationFromSourceZRot
0021|GEMS_RELA_01|54|SH|3|ImagePosition
0021|GEMS_RELA_01|55|SH|6|ImageOrientation
0021|GEMS_RELA_01|56|SL|1|IntegerSlop
0021|GEMS_RELA_01|57|SL|1|IntegerSlop
0021|GEMS_RELA_01|58|SL|1|IntegerSlop
0021|GEMS_RELA_01|59|SL|1|IntegerSlop
0021|GEMS_RELA_01|5a|SL|1|IntegerSlop
0021|GEMS_RELA_01|5b|DS|1|FloatSlop
0021|GEMS_RELA_01|5c|DS|1|FloatSlop
0021|GEMS_RELA_01|5d|DS|1|FloatSlop
0021|GEMS_RELA_01|5e|DS|1|FloatSlop
0021|GEMS_RELA_01|5f|DS|1|FloatSlop
0021|GEMS_RELA_01|81|DS|1|AutoWindowLevelAlpha
0021|GEMS_RELA_01|83|DS|1|AutoWindowLevelWindow
0021|GEMS_RELA_01|84|DS|1|AutoWindowLevelLevel
0043|GEMS_PARM_01|36|UL|1|UserFillMapMSW
0043|GEMS_PARM_01|37|UL|1|UserFillMapLSW
0043|GEMS_PARM_01|38|FL|24|User25ToUser48
0043|GEMS_PARM_01|39|IS|4|SlopInteger6ToSlopInteger9
0043|GEMS_PARM_01|40|FL|4|TriggerOnPosition
0043|GEMS_PARM_01|41|FL|4|DegreeOfRotation
0043|GEMS_PARM_01|42|SL|4|DASTriggerSource
0043|GEMS_PARM_01|43|SL|4|DASFpaGain
0043|GEMS_PARM_01|44|SL|4|DASOutputSource
0043|GEMS_PARM_01|45|SL|4|DASAdInput
0043|GEMS_PARM_01|46|SL|4|DASCalMode
0043|GEMS_PARM_01|47|SL|4|DASCalFrequency
0043|GEMS_PARM_01|48|SL|4|DASRegXm
0043|GEMS_PARM_01|49|SL|4|DASAutoZero
0043|GEMS_PARM_01|4a|SS|4|StartingChannelOfView
0043|GEMS_PARM_01|4b|SL|4|DASXmPattern
0043|GEMS_PARM_01|4c|SS|4|TGGCTriggerMode
0043|GEMS_PARM_01|4d|FL|4|StartScanToXrayOnDelay
0043|GEMS_PARM_01|60|IS|8|Unknown
0043|GEMS_PARM_01|61|UI|1|Unknown
0043|GEMS_PARM_01|62|SH|1|Unknown
0043|GEMS_PARM_01|6f|DS|3|Unknown
0045|GEMS_SENO_02|04|CS|1|AES
0045|GEMS_SENO_02|06|DS|1|Angulation
0045|GEMS_SENO_02|09|DS|1|RealMagnificationFactor
0045|GEMS_SENO_02|0b|CS|1|SenographType
0045|GEMS_SENO_02|0c|DS|1|IntegrationTime
0045|GEMS_SENO_02|0d|DS|1|ROIOriginXY
0045|GEMS_SENO_02|11|DS|2|ReceptorSizeCmXY
0045|GEMS_SENO_02|12|IS|2|ReceptorSizePixelsXY
0045|GEMS_SENO_02|13|ST|1|Screen
0045|GEMS_SENO_02|14|DS|1|PixelPitchMicrons
0045|GEMS_SENO_02|15|IS|1|PixelDepthBits
0045|GEMS_SENO_02|16|IS|2|BinningFactorXY
0045|GEMS_SENO_02|1B|CS|1|ClinicalView
0045|GEMS_SENO_02|1D|DS|1|MeanOfRawGrayLevels
0045|GEMS_SENO_02|1E|DS|1|MeanOfOffsetGrayLevels
0045|GEMS_SENO_02|1F|DS|1|MeanOfCorrectedGrayLevels
0045|GEMS_SENO_02|20|DS|1|MeanOfRegionGrayLevels
0045|GEMS_SENO_02|21|DS|1|MeanOfLogRegionGrayLevels
0045|GEMS_SENO_02|22|DS|1|StandardDeviationOfRawGrayLevels
0045|GEMS_SENO_02|23|DS|1|StandardDeviationOfCorrectedGrayLevels
0045|GEMS_SENO_02|24|DS|1|StandardDeviationOfRegionGrayLevels
0045|GEMS_SENO_02|25|DS|1|StandardDeviationOfLogRegionGrayLevels
0045|GEMS_SENO_02|26|OB|1|MAOBuffer
0045|GEMS_SENO_02|27|IS|1|SetNumber
0045|GEMS_SENO_02|28|CS|1|WindowingType
0045|GEMS_SENO_02|29|DS|1-n|WindowingParameters
0045|GEMS_SENO_02|2a|IS|1|CrosshairCursorXCoordinates
0045|GEMS_SENO_02|2b|IS|1|CrosshairCursorYCoordinates
0045|GEMS_SENO_02|39|US|1|VignetteRows
0045|GEMS_SENO_02|3a|US|1|VignetteColumns
0045|GEMS_SENO_02|3b|US|1|VignetteBitsAllocated
0045|GEMS_SENO_02|3c|US|1|VignetteBitsStored
0045|GEMS_SENO_02|3d|US|1|VignetteHighBit
0045|GEMS_SENO_02|3e|US|1|VignettePixelRepresentation
0045|GEMS_SENO_02|3f|OB|1|VignettePixelData
0033|GEMS_YMHD_01|05|UN|1|Unknown
0033|GEMS_YMHD_01|06|UN|1|Unknown
0019|GE_GENESIS_REV3.0|39|SS|1|AxialType
0019|SVISION|78|DS|1|FilterThickness1
0021|GEMS_RELA_01|91|SS|1|BiopsyPosition
0021|GEMS_RELA_01|93|FL|1|BiopsyRefLocation
0023|GEMS_STDY_01|01|SL|1|NumberOfSeriesInStudy
0023|GEMS_STDY_01|02|SL|1|NumberOfUnarchivedSeries
0023|GEMS_STDY_01|10|SS|1|ReferenceImageField
0023|GEMS_STDY_01|50|SS|1|SummaryImage
0023|GEMS_STDY_01|70|FD|1|StartTimeSecsInFirstAxial
0023|GEMS_STDY_01|74|SL|1|NumberOfUpdatesToHeader
0023|GEMS_STDY_01|7d|SS|1|IndicatesIfStudyHasCompleteInfo
0025|GEMS_SERS_01|06|SS|1|LastPulseSequenceUsed
0025|GEMS_SERS_01|07|SL|1|ImagesInSeries
0025|GEMS_SERS_01|10|SL|1|LandmarkCounter
0025|GEMS_SERS_01|11|SS|1|NumberOfAcquisitions
0025|GEMS_SERS_01|14|SL|1|IndicatesNumberOfUpdatesToHeader
0025|GEMS_SERS_01|17|SL|1|SeriesCompleteFlag
0025|GEMS_SERS_01|18|SL|1|NumberOfImagesArchived
0025|GEMS_SERS_01|19|SL|1|LastImageNumberUsed
0025|GEMS_SERS_01|1a|SH|1|PrimaryReceiverSuiteAndHost
0019|GE_GENESIS_REV3.0|8f|SS|1|SwapPhaseFrequency
0019|GE_GENESIS_REV3.0|9c|SS|1|PulseSequenceName
0019|GE_GENESIS_REV3.0|9f|SS|1|CoilType
0019|GE_GENESIS_REV3.0|a4|SS|1|SATFatWaterBone
0019|GE_GENESIS_REV3.0|c0|SS|1|BitmapOfSATSelections
0019|GE_GENESIS_REV3.0|c1|SS|1|SurfaceCoilIntensityCorrectionFlag
0019|GE_GENESIS_REV3.0|cb|SS|1|PhaseContrastFlowAxis
0019|GE_GENESIS_REV3.0|cc|SS|1|PhaseContrastVelocityEncoding
0019|GE_GENESIS_REV3.0|d5|SS|1|FractionalEcho
0019|GE_GENESIS_REV3.0|d8|SS|1|VariableEchoFlag
0019|GE_GENESIS_REV3.0|d9|DS|1|ConcatenatedSat
0019|GE_GENESIS_REV3.0|f2|SS|1|NumberOfPhases
0043|GE_GENESIS_REV3.0|1e|DS|1|DeltaStartTime
0043|GE_GENESIS_REV3.0|27|SH|1|ScanPitchRatio
0029|INTELERAD MEDICAL SYSTEMS|01|FD|1|ImageCompressionFraction
0029|INTELERAD MEDICAL SYSTEMS|02|FD|1|ImageQuality
0029|INTELERAD MEDICAL SYSTEMS|03|FD|1|ImageBytesTransferred
0029|INTELERAD MEDICAL SYSTEMS|10|SH|1|J2cParameterType
0029|INTELERAD MEDICAL SYSTEMS|11|US|1|J2cPixelRepresentation
0029|INTELERAD MEDICAL SYSTEMS|12|US|1|J2cBitsAllocated
0029|INTELERAD MEDICAL SYSTEMS|13|US|1|J2cPixelShiftValue
0029|INTELERAD MEDICAL SYSTEMS|14|US|1|J2cPlanarConfiguration
0029|INTELERAD MEDICAL SYSTEMS|15|DS|1|J2cRescaleIntercept
0029|INTELERAD MEDICAL SYSTEMS|20|LO|1|PixelDataMD5SumPerFrame
0029|INTELERAD MEDICAL SYSTEMS|21|US|1|HistogramPercentileLabels
0029|INTELERAD MEDICAL SYSTEMS|22|FD|1|HistogramPercentileValues
3f01|INTELERAD MEDICAL SYSTEMS|01|LO|1|InstitutionCode
3f01|INTELERAD MEDICAL SYSTEMS|02|LO|1|RoutedTransferAE
3f01|INTELERAD MEDICAL SYSTEMS|03|LO|1|SourceAE
3f01|INTELERAD MEDICAL SYSTEMS|04|SH|1|DeferredValidation
3f01|INTELERAD MEDICAL SYSTEMS|05|LO|1|SeriesOwner
3f01|INTELERAD MEDICAL SYSTEMS|06|LO|1|OrderGroupNumber
3f01|INTELERAD MEDICAL SYSTEMS|07|SH|1|StrippedPixelData
3f01|INTELERAD MEDICAL SYSTEMS|08|SH|1|PendingMoveRequest
0041|INTEGRIS 1.0|20|FL|1|AccumulatedFluoroscopyDose
0041|INTEGRIS 1.0|30|FL|1|AccumulatedExposureDose
0041|INTEGRIS 1.0|40|FL|1|TotalDose
0041|INTEGRIS 1.0|41|FL|1|TotalNumberOfFrames
0041|INTEGRIS 1.0|50|SQ|1|ExposureInformationSequence
0009|INTEGRIS 1.0|08|CS|1-n|ExposureChannel
0009|INTEGRIS 1.0|32|TM|1|ExposureStartTime
0019|INTEGRIS 1.0|00|LO|1|APRName
0019|INTEGRIS 1.0|40|DS|1|FrameRate
0021|INTEGRIS 1.0|12|IS|1|ExposureNumber
0029|INTEGRIS 1.0|08|IS|1|NumberOfExposureResults
0029|ISG shadow|70|IS|1|Unknown
0029|ISG shadow|80|IS|1|Unknown
0029|ISG shadow|90|IS|1|Unknown
0009|ISI|01|UN|1|SIENETGeneralPurposeIMGEF
0009|MERGE TECHNOLOGIES, INC.|00|OB|1|Unknown
0029|OCULUS Optikgeraete GmbH|1010|OB|1|OriginalMeasuringData
0019|SVISION|79|DS|1|FilterThickness2
0029|OCULUS Optikgeraete GmbH|1012|UL|1|OriginalMeasuringDataLength
0029|OCULUS Optikgeraete GmbH|1020|OB|1|OriginalMeasuringRawData
0029|OCULUS Optikgeraete GmbH|1022|UL|1|OriginalMeasuringRawDataLength
0041|PAPYRUS 3.0|00|LT|1|PapyrusComments
0041|PAPYRUS 3.0|10|SQ|1|PointerSequence
0041|PAPYRUS 3.0|11|UL|1|ImagePointer
0041|PAPYRUS 3.0|12|UL|1|PixelOffset
0041|PAPYRUS 3.0|13|SQ|1|ImageIdentifierSequence
0041|PAPYRUS 3.0|14|SQ|1|ExternalFileReferenceSequence
0041|PAPYRUS 3.0|15|US|1|NumberOfImages
0041|PAPYRUS 3.0|21|UI|1|ReferencedSOPClassUID
0041|PAPYRUS 3.0|22|UI|1|ReferencedSOPInstanceUID
0041|PAPYRUS 3.0|31|LT|1|ReferencedFileName
0041|PAPYRUS 3.0|32|LT|1-n|ReferencedFilePath
0041|PAPYRUS 3.0|41|UI|1|ReferencedImageSOPClassUID
0041|PAPYRUS 3.0|42|UI|1|ReferencedImageSOPInstanceUID
0041|PAPYRUS 3.0|50|SQ|1|ImageSequence
0009|PAPYRUS|00|LT|1|OriginalFileName
0009|PAPYRUS|10|LT|1|OriginalFileLocation
0009|PAPYRUS|18|LT|1|DataSetIdentifier
0041|PAPYRUS|00|LT|1-n|PapyrusComments
0041|PAPYRUS|10|US|1|FolderType
0041|PAPYRUS|11|LT|1|PatientFolderDataSetID
0041|PAPYRUS|20|LT|1|FolderName
0041|PAPYRUS|30|DA|1|CreationDate
0041|PAPYRUS|32|TM|1|CreationTime
0041|PAPYRUS|34|DA|1|ModifiedDate
0041|PAPYRUS|36|TM|1|ModifiedTime
0041|PAPYRUS|40|LT|1-n|OwnerName
0041|PAPYRUS|50|LT|1|FolderStatus
0041|PAPYRUS|60|UL|1|NumberOfImages
0041|PAPYRUS|62|UL|1|NumberOfOther
0041|PAPYRUS|a0|LT|1-n|ExternalFolderElementDSID
0041|PAPYRUS|a1|US|1-n|ExternalFolderElementDataSetType
0041|PAPYRUS|a2|LT|1-n|ExternalFolderElementFileLocation
0041|PAPYRUS|a3|UL|1-n|ExternalFolderElementLength
0041|PAPYRUS|b0|LT|1-n|InternalFolderElementDSID
0041|PAPYRUS|b1|US|1-n|InternalFolderElementDataSetType
0041|PAPYRUS|b2|UL|1-n|InternalOffsetToDataSet
0041|PAPYRUS|b3|UL|1-n|InternalOffsetToImage
2001|Philips Imaging DD 001|17|SL|1|NumberOfPhasesMR
2001|Philips Imaging DD 001|18|SL|1|NumberOfSlicesMR
2001|Philips Imaging DD 001|3f|CS|1|ZoomMode
2001|Philips Imaging DD 001|62|CS|1|SeriesCommitted
2001|PHILIPS IMAGING DD 001|01|FL|1|ChemicalShift
2001|PHILIPS IMAGING DD 001|02|IS|1|ChemicalShiftNumberMR
2001|PHILIPS IMAGING DD 001|03|FL|1|DiffusionB-Factor
2001|PHILIPS IMAGING DD 001|04|CS|1|DiffusionDirection
2001|PHILIPS IMAGING DD 001|06|CS|1|ImageEnhanced
2001|PHILIPS IMAGING DD 001|07|CS|1|ImageTypeEDES
2001|PHILIPS IMAGING DD 001|08|IS|1|PhaseNumber
2001|PHILIPS IMAGING DD 001|0a|IS|1|SliceNumberMR
2001|PHILIPS IMAGING DD 001|0b|CS|1|SliceOrientation
2001|PHILIPS IMAGING DD 001|11|FL|1|DiffusionEchoTime
2001|PHILIPS IMAGING DD 001|12|CS|1|DynamicSeries
2001|PHILIPS IMAGING DD 001|13|SL|1|EPIFactor
2001|PHILIPS IMAGING DD 001|14|SL|1|NumberOfEchoes
2001|PHILIPS IMAGING DD 001|15|SS|1|NumberOfLocations
2001|PHILIPS IMAGING DD 001|16|SS|1|NumberOfPCDirections
2001|PHILIPS IMAGING DD 001|17|SL|1|NumberOfPhasesMR
2001|PHILIPS IMAGING DD 001|18|SL|1|NumberOfSlicesMR
2001|PHILIPS IMAGING DD 001|19|CS|1|PartialMatrixScanned
2001|PHILIPS IMAGING DD 001|1a|FL|1-n|PCVelocity
2001|PHILIPS IMAGING DD 001|1b|FL|1|PrepulseDelay
2001|PHILIPS IMAGING DD 001|1c|CS|1|PrepulseType
2001|PHILIPS IMAGING DD 001|1d|IS|1|ReconstructionNumberMR
2001|PHILIPS IMAGING DD 001|1f|CS|1|RespirationSync
2001|PHILIPS IMAGING DD 001|21|CS|1|SPIR
2001|PHILIPS IMAGING DD 001|22|FL|1|WaterFatShift
2001|PHILIPS IMAGING DD 001|23|DS|1|FlipAnglePhilips
2001|Philips Imaging DD 001|1a|FL|1-n|PCVelocity
2001|PHILIPS IMAGING DD 001|25|SH|1|EchoTimeDisplayMR
2001|PHILIPS IMAGING DD 001|2d|SS|1|StackNumberOfSlices
2001|PHILIPS IMAGING DD 001|32|FL|1|StackRadialAngle
2001|PHILIPS IMAGING DD 001|33|CS|1|StackRadialAxis
2001|PHILIPS IMAGING DD 001|35|SS|1|StackSliceNumber
2001|PHILIPS IMAGING DD 001|36|CS|1|StackType
2001|PHILIPS IMAGING DD 001|3f|CS|1|ZoomMode
2001|PHILIPS IMAGING DD 001|5f|SQ|1-n|StackSequence
2001|PHILIPS IMAGING DD 001|60|SL|1|NumberOfStacks
2001|PHILIPS IMAGING DD 001|61|CS|1|SeriesTransmitted
2001|PHILIPS IMAGING DD 001|62|CS|1|SeriesCommitted
2001|PHILIPS IMAGING DD 001|63|CS|1|ExaminationSource
2001|PHILIPS IMAGING DD 001|7b|IS|1|AcquisitionNumber
2001|PHILIPS IMAGING DD 001|81|IS|1|NumberOfDynamicScans
2005|Philips MR Imaging DD 001|05|CS|1|SynergyReconstructionType
2005|Philips MR Imaging DD 001|1e|SH|1|MIPProtocol
2005|Philips MR Imaging DD 001|1f|SH|1|MPRProtocol
2005|Philips MR Imaging DD 001|2d|SS|1|NumberOfStackSlices
2005|Philips MR Imaging DD 001|32|FL|1|StackRadialAngle
2005|Philips MR Imaging DD 001|33|CS|1|StackRadialAxis
2005|Philips MR Imaging DD 001|35|SS|1|StackSliceNumber
2005|Philips MR Imaging DD 001|36|CS|1|StackType
2005|Philips MR Imaging DD 001|5f|SQ|1|StackSequence
2005|Philips MR Imaging DD 001|83|SQ|1|Unknown
2005|Philips MR Imaging DD 005|02|SQ|1|Unknown
2005|PHILIPS MR IMAGING DD 001|05|CS|1|SynergyReconstructionType
2005|PHILIPS MR IMAGING DD 001|1e|SH|1|MIPProtocol
2005|PHILIPS MR IMAGING DD 001|1f|SH|1|MPRProtocol
2005|PHILIPS MR IMAGING DD 001|20|SL|1|NumberOfChemicalShifts
2005|PHILIPS MR IMAGING DD 001|2d|SS|1|NumberOfStackSlices
2005|PHILIPS MR IMAGING DD 001|32|FL|1|StackRadialAngle
2005|PHILIPS MR IMAGING DD 001|33|CS|1|StackRadialAxis
2005|PHILIPS MR IMAGING DD 001|35|SS|1|StackSliceNumber
2005|PHILIPS MR IMAGING DD 001|36|CS|1|StackType
2005|PHILIPS MR IMAGING DD 001|a1|CS|1|SyncraScanType
2005|PHILIPS MR IMAGING DD 001|5f|SQ|1|StackSequence
2005|PHILIPS MR IMAGING DD 001|83|SQ|1|Unknown
0019|PHILIPS MR R5.5/PART|1000|DS|1|FieldOfView
0019|PHILIPS MR R5.6/PART|1000|DS|1|FieldOfView
0019|PHILIPS MR SPECTRO;1|01|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|02|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|03|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|04|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|05|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|06|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|07|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|08|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|09|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|10|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|12|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|13|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|14|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|15|US|1-n|Unknown
0019|PHILIPS MR SPECTRO;1|16|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|17|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|18|UN|1|Unknown
0019|PHILIPS MR SPECTRO;1|20|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|21|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|22|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|23|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|24|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|25|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|26|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|27|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|28|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|29|IS|1-n|Unknown
0019|PHILIPS MR SPECTRO;1|31|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|32|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|41|LT|1|Unknown
0019|PHILIPS MR SPECTRO;1|42|IS|2|Unknown
0019|PHILIPS MR SPECTRO;1|43|IS|2|Unknown
0019|PHILIPS MR SPECTRO;1|45|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|46|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|47|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|48|IS|1|Unknown
0019|PHILIPS MR SPECTRO;1|49|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|50|UN|1|Unknown
0019|PHILIPS MR SPECTRO;1|60|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|61|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|70|UN|1|Unknown
0019|PHILIPS MR SPECTRO;1|71|IS|1-n|Unknown
0019|PHILIPS MR SPECTRO;1|72|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|73|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|74|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|76|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|77|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|78|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|79|US|1|Unknown
0019|PHILIPS MR SPECTRO;1|80|IS|1|Unknown
0009|PHILIPS MR|10|LO|1|SPIRelease
0009|PHILIPS MR|12|LO|1|Unknown
0019|PHILIPS MR/LAST|09|DS|1|MainMagneticField
0019|PHILIPS MR/LAST|0e|IS|1|FlowCompensation
0019|PHILIPS MR/LAST|b1|IS|1|MinimumRRInterval
0019|PHILIPS MR/LAST|b2|IS|1|MaximumRRInterval
0019|PHILIPS MR/LAST|b3|IS|1|NumberOfRejections
0019|PHILIPS MR/LAST|b4|IS|1-n|NumberOfRRIntervals
0019|PHILIPS MR/LAST|b5|IS|1|ArrhythmiaRejection
0019|PHILIPS MR/LAST|c0|DS|1-n|Unknown
0019|PHILIPS MR/LAST|c6|IS|1|CycledMultipleSlice
0019|PHILIPS MR/LAST|ce|IS|1|REST
0019|PHILIPS MR/LAST|d5|DS|1|Unknown
0019|PHILIPS MR/LAST|d6|IS|1|FourierInterpolation
0019|PHILIPS MR/LAST|d9|IS|1-n|Unknown
0019|PHILIPS MR/LAST|e0|IS|1|Prepulse
0019|PHILIPS MR/LAST|e1|DS|1|PrepulseDelay
0019|PHILIPS MR/LAST|e2|IS|1|Unknown
0019|PHILIPS MR/LAST|e3|DS|1|Unknown
0019|PHILIPS MR/LAST|f0|LT|1|WSProtocolString1
0019|PHILIPS MR/LAST|f1|LT|1|WSProtocolString2
0019|PHILIPS MR/LAST|f2|LT|1|WSProtocolString3
0019|PHILIPS MR/LAST|f3|LT|1|WSProtocolString4
0021|PHILIPS MR/LAST|00|IS|1|Unknown
0021|PHILIPS MR/LAST|10|IS|1|Unknown
0021|PHILIPS MR/LAST|20|IS|1|Unknown
0021|PHILIPS MR/LAST|21|DS|1|SliceGap
0021|PHILIPS MR/LAST|22|DS|1|StackRadialAngle
0027|PHILIPS MR/LAST|00|US|1|Unknown
0027|PHILIPS MR/LAST|11|US|1-n|Unknown
0027|PHILIPS MR/LAST|12|DS|1-n|Unknown
0027|PHILIPS MR/LAST|13|DS|1-n|Unknown
0027|PHILIPS MR/LAST|14|DS|1-n|Unknown
0027|PHILIPS MR/LAST|15|DS|1-n|Unknown
0027|PHILIPS MR/LAST|16|LO|1|Unknown
0029|PHILIPS MR/LAST|10|DS|1|FPMin
0029|PHILIPS MR/LAST|20|DS|1|FPMax
0029|PHILIPS MR/LAST|30|DS|1|ScaledMinimum
0029|PHILIPS MR/LAST|40|DS|1|ScaledMaximum
0029|PHILIPS MR/LAST|50|DS|1|WindowMinimum
0029|PHILIPS MR/LAST|60|DS|1|WindowMaximum
0029|PHILIPS MR/LAST|61|IS|1|Unknown
0029|PHILIPS MR/LAST|70|DS|1|Unknown
0029|PHILIPS MR/LAST|71|DS|1|Unknown
0029|PHILIPS MR/LAST|72|IS|1|Unknown
0029|PHILIPS MR/LAST|80|IS|1|ViewCenter
0029|PHILIPS MR/LAST|81|IS|1|ViewSize
0029|PHILIPS MR/LAST|82|IS|1|ViewZoom
0029|PHILIPS MR/LAST|83|IS|1|ViewTransform
6001|PHILIPS MR/LAST|00|LT|1|Unknown
0019|PHILIPS MR/PART|1000|DS|1|FieldOfView
0019|PHILIPS MR/PART|1005|DS|1|CCAngulation
0019|PHILIPS MR/PART|1006|DS|1|APAngulation
0019|PHILIPS MR/PART|1007|DS|1|LRAngulation
0019|PHILIPS MR/PART|1008|IS|1|PatientPosition
0019|PHILIPS MR/PART|1009|IS|1|PatientOrientation
0019|PHILIPS MR/PART|100a|IS|1|SliceOrientation
0019|PHILIPS MR/PART|100b|DS|1|LROffcenter
0019|PHILIPS MR/PART|100c|DS|1|CCOffcenter
0019|PHILIPS MR/PART|100d|DS|1|APOffcenter
0019|PHILIPS MR/PART|100e|DS|1|Unknown
0019|PHILIPS MR/PART|100f|IS|1|NumberOfSlices
0019|PHILIPS MR/PART|1010|DS|1|SliceFactor
0019|PHILIPS MR/PART|1011|DS|1-n|EchoTimes
0019|PHILIPS MR/PART|1015|IS|1|DynamicStudy
0019|PHILIPS MR/PART|1018|DS|1|HeartbeatInterval
0019|PHILIPS MR/PART|1019|DS|1|RepetitionTimeFFE
0019|PHILIPS MR/PART|101a|DS|1|FFEFlipAngle
0019|PHILIPS MR/PART|101b|IS|1|NumberOfScans
0019|PHILIPS MR/PART|1021|DS|1-n|Unknown
0019|PHILIPS MR/PART|1022|DS|1|DynamicScanTimeBegin
0019|PHILIPS MR/PART|1024|IS|1|Unknown
0019|PHILIPS MR/PART|1064|DS|1|RepetitionTimeSE
0019|PHILIPS MR/PART|1065|DS|1|RepetitionTimeIR
0019|PHILIPS MR/PART|1069|IS|1|NumberOfPhases
0019|PHILIPS MR/PART|106a|IS|1|CardiacFrequency
0019|PHILIPS MR/PART|106b|DS|1|InversionDelay
0019|PHILIPS MR/PART|106c|DS|1|GateDelay
0019|PHILIPS MR/PART|106d|DS|1|GateWidth
0019|PHILIPS MR/PART|106e|DS|1|TriggerDelayTime
0019|PHILIPS MR/PART|1080|IS|1|NumberOfChemicalShifts
0019|PHILIPS MR/PART|1081|DS|1|ChemicalShift
0019|PHILIPS MR/PART|1084|IS|1|NumberOfRows
0019|PHILIPS MR/PART|1085|IS|1|NumberOfSamples
0019|PHILIPS MR/PART|1094|LO|1|MagnetizationTransferContrast
0019|PHILIPS MR/PART|1095|LO|1|SpectralPresaturationWithInversionRecovery
0019|PHILIPS MR/PART|1096|IS|1|Unknown
0019|PHILIPS MR/PART|1097|LO|1|Unknown
0019|PHILIPS MR/PART|10a0|IS|1|Unknown
0019|PHILIPS MR/PART|10a1|DS|1|Unknown
0019|PHILIPS MR/PART|10a3|DS|1|Unknown
0019|PHILIPS MR/PART|10a4|CS|1|Unknown
0019|PHILIPS MR/PART|10c8|IS|1|Unknown
0019|PHILIPS MR/PART|10c9|IS|1|FoldoverDirectionTransverse
0019|PHILIPS MR/PART|10ca|IS|1|FoldoverDirectionSagittal
0019|PHILIPS MR/PART|10cb|IS|1|FoldoverDirectionCoronal
0019|PHILIPS MR/PART|10cc|IS|1|Unknown
0019|PHILIPS MR/PART|10cd|IS|1|Unknown
0019|PHILIPS MR/PART|10ce|IS|1|Unknown
0019|PHILIPS MR/PART|10cf|IS|1|NumberOfEchoes
0019|PHILIPS MR/PART|10d0|IS|1|ScanResolution
0019|PHILIPS MR/PART|10d2|LO|2|WaterFatShift
0019|PHILIPS MR/PART|10d4|IS|1|ArtifactReduction
0019|PHILIPS MR/PART|10d5|IS|1|Unknown
0019|PHILIPS MR/PART|10d6|IS|1|Unknown
0019|PHILIPS MR/PART|10d7|DS|1|ScanPercentage
0019|PHILIPS MR/PART|10d8|IS|1|Halfscan
0019|PHILIPS MR/PART|10d9|IS|1|EPIFactor
0019|PHILIPS MR/PART|10da|IS|1|TurboFactor
0019|PHILIPS MR/PART|10db|IS|1|Unknown
0019|PHILIPS MR/PART|10e0|IS|1|PercentageOfScanCompleted
0019|PHILIPS MR/PART|10e1|IS|1|Unknown
0019|PHILIPS MR/PART|1100|IS|1|NumberOfStacks
0019|PHILIPS MR/PART|1101|IS|1-n|StackType
0019|PHILIPS MR/PART|1102|IS|1-n|Unknown
0019|PHILIPS MR/PART|110b|DS|1|LROffcenter
0019|PHILIPS MR/PART|110c|DS|1|CCOffcenter
0019|PHILIPS MR/PART|110d|DS|1|APOffcenter
0019|PHILIPS MR/PART|1145|IS|1|ReconstructionResolution
0019|PHILIPS MR/PART|11fc|IS|1|ResonanceFrequency
0019|PHILIPS MR/PART|12c0|DS|1|TriggerDelayTimes
0019|PHILIPS MR/PART|12e0|IS|1|PrepulseType
0019|PHILIPS MR/PART|12e1|DS|1|PrepulseDelay
0019|PHILIPS MR/PART|12e3|DS|1|PhaseContrastVelocity
0021|PHILIPS MR/PART|1000|IS|1|ReconstructionNumber
0021|PHILIPS MR/PART|1010|IS|1|ImageType
0021|PHILIPS MR/PART|1020|IS|1|SliceNumber
0021|PHILIPS MR/PART|1030|IS|1|EchoNumber
0021|PHILIPS MR/PART|1031|DS|1|PatientReferenceID
0021|PHILIPS MR/PART|1035|IS|1|ChemicalShiftNumber
0021|PHILIPS MR/PART|1040|IS|1|PhaseNumber
0021|PHILIPS MR/PART|1050|IS|1|DynamicScanNumber
0021|PHILIPS MR/PART|1060|IS|1|NumberOfRowsInObject
0021|PHILIPS MR/PART|1061|IS|1-n|RowNumber
0021|PHILIPS MR/PART|1062|IS|1-n|Unknown
0021|PHILIPS MR/PART|1100|DA|1|ScanDate
0021|PHILIPS MR/PART|1110|TM|1|ScanTime
0021|PHILIPS MR/PART|1221|IS|1|SliceGap
0029|PHILIPS MR/PART|00|DS|2|Unknown
0029|PHILIPS MR/PART|04|US|1|Unknown
0029|PHILIPS MR/PART|10|DS|1|Unknown
0029|PHILIPS MR/PART|11|DS|1|Unknown
0029|PHILIPS MR/PART|20|LO|1|Unknown
0029|PHILIPS MR/PART|31|DS|2|Unknown
0029|PHILIPS MR/PART|32|DS|2|Unknown
0029|PHILIPS MR/PART|c3|IS|1|ScanResolution
0029|PHILIPS MR/PART|c4|IS|1|FieldOfView
0029|PHILIPS MR/PART|d5|LT|1|SliceThickness
0019|PHILIPS-MR-1|11|IS|1|ChemicalShiftNumber
0019|PHILIPS-MR-1|12|IS|1|PhaseNumber
0021|PHILIPS-MR-1|01|IS|1|ReconstructionNumber
0021|PHILIPS-MR-1|02|IS|1|SliceNumber
7001|Picker NM Private Group|01|UI|1|Unknown
7001|Picker NM Private Group|02|OB|1|Unknown
0019|SIEMENS CM VA0  ACQU|10|LT|1|ParameterFileName
0019|SIEMENS CM VA0  ACQU|11|LO|1|SequenceFileName
0019|SIEMENS CM VA0  ACQU|12|LT|1|SequenceFileOwner
0019|SIEMENS CM VA0  ACQU|13|LT|1|SequenceDescription
0019|SIEMENS CM VA0  ACQU|14|LT|1|EPIFileName
0009|SIEMENS CM VA0  CMS|00|DS|1|NumberOfMeasurements
0009|SIEMENS CM VA0  CMS|10|LT|1|StorageMode
0009|SIEMENS CM VA0  CMS|12|UL|1|EvaluationMaskImage
0009|SIEMENS CM VA0  CMS|26|DA|1|LastMoveDate
0009|SIEMENS CM VA0  CMS|27|TM|1|LastMoveTime
0011|SIEMENS CM VA0  CMS|0a|LT|1|Unknown
0011|SIEMENS CM VA0  CMS|10|DA|1|RegistrationDate
0011|SIEMENS CM VA0  CMS|11|TM|1|RegistrationTime
0011|SIEMENS CM VA0  CMS|22|LT|1|Unknown
0011|SIEMENS CM VA0  CMS|23|DS|1|UsedPatientWeight
0011|SIEMENS CM VA0  CMS|40|IS|1|OrganCode
0013|SIEMENS CM VA0  CMS|00|LT|1|ModifyingPhysician
0013|SIEMENS CM VA0  CMS|10|DA|1|ModificationDate
0013|SIEMENS CM VA0  CMS|12|TM|1|ModificationTime
0013|SIEMENS CM VA0  CMS|20|LO|1|PatientName
0013|SIEMENS CM VA0  CMS|22|LO|1|PatientId
0013|SIEMENS CM VA0  CMS|30|DA|1|PatientBirthdate
0013|SIEMENS CM VA0  CMS|31|DS|1|PatientWeight
0013|SIEMENS CM VA0  CMS|32|LT|1|PatientsMaidenName
0013|SIEMENS CM VA0  CMS|33|LT|1|ReferringPhysician
0013|SIEMENS CM VA0  CMS|34|LT|1|AdmittingDiagnosis
0013|SIEMENS CM VA0  CMS|35|LO|1|PatientSex
0013|SIEMENS CM VA0  CMS|40|LO|1|ProcedureDescription
0013|SIEMENS CM VA0  CMS|42|LO|1|RestDirection
0013|SIEMENS CM VA0  CMS|44|LO|1|PatientPosition
0013|SIEMENS CM VA0  CMS|46|LT|1|ViewDirection
0013|SIEMENS CM VA0  CMS|50|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|51|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|52|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|53|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|54|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|55|LT|1|Unknown
0013|SIEMENS CM VA0  CMS|56|LT|1|Unknown
0019|SIEMENS CM VA0  CMS|10|DS|1|NetFrequency
0019|SIEMENS CM VA0  CMS|20|LT|1|MeasurementMode
0019|SIEMENS CM VA0  CMS|30|LT|1|CalculationMode
0019|SIEMENS CM VA0  CMS|50|IS|1|NoiseLevel
0019|SIEMENS CM VA0  CMS|60|IS|1|NumberOfDataBytes
0021|SIEMENS CM VA0  CMS|20|DS|2|FoV
0021|SIEMENS CM VA0  CMS|22|DS|1|ImageMagnificationFactor
0021|SIEMENS CM VA0  CMS|24|DS|2|ImageScrollOffset
0021|SIEMENS CM VA0  CMS|26|IS|1|ImagePixelOffset
0021|SIEMENS CM VA0  CMS|30|LT|1|ViewDirection
0021|SIEMENS CM VA0  CMS|32|CS|1|PatientRestDirection
0021|SIEMENS CM VA0  CMS|60|DS|3|ImagePosition
0021|SIEMENS CM VA0  CMS|61|DS|3|ImageNormal
0021|SIEMENS CM VA0  CMS|63|DS|1|ImageDistance
0021|SIEMENS CM VA0  CMS|65|US|1|ImagePositioningHistoryMask
0021|SIEMENS CM VA0  CMS|6a|DS|3|ImageRow
0021|SIEMENS CM VA0  CMS|6b|DS|3|ImageColumn
0021|SIEMENS CM VA0  CMS|70|LT|3|PatientOrientationSet1
0021|SIEMENS CM VA0  CMS|71|LT|3|PatientOrientationSet2
0021|SIEMENS CM VA0  CMS|80|LT|1|StudyName
0021|SIEMENS CM VA0  CMS|82|LT|3|StudyType
0029|SIEMENS CM VA0  CMS|10|LT|1|WindowStyle
0029|SIEMENS CM VA0  CMS|11|LT|1|Unknown
0029|SIEMENS CM VA0  CMS|13|LT|1|Unknown
0029|SIEMENS CM VA0  CMS|20|LT|3|PixelQualityCode
0029|SIEMENS CM VA0  CMS|22|IS|3|PixelQualityValue
0029|SIEMENS CM VA0  CMS|50|LT|1|ArchiveCode
0029|SIEMENS CM VA0  CMS|51|LT|1|ExposureCode
0029|SIEMENS CM VA0  CMS|52|LT|1|SortCode
0029|SIEMENS CM VA0  CMS|53|LT|1|Unknown
0029|SIEMENS CM VA0  CMS|60|LT|1|Splash
0051|SIEMENS CM VA0  CMS|10|LT|1-n|ImageText
6021|SIEMENS CM VA0  CMS|00|LT|1|ImageGraphicsFormatCode
6021|SIEMENS CM VA0  CMS|10|LT|1|ImageGraphics
7fe1|SIEMENS CM VA0  CMS|00|OB|1-n|BinaryData
0009|SIEMENS CM VA0  LAB|10|LT|1|GeneratorIdentificationLabel
0009|SIEMENS CM VA0  LAB|11|LT|1|GantryIdentificationLabel
0009|SIEMENS CM VA0  LAB|12|LT|1|X-RayTubeIdentificationLabel
0019|SVISION|80|IS|1|BuckyFormat
0009|SIEMENS CM VA0  LAB|13|LT|1|DetectorIdentificationLabel
0009|SIEMENS CM VA0  LAB|14|LT|1|DASIdentificationLabel
0009|SIEMENS CM VA0  LAB|15|LT|1|SMIIdentificationLabel
0009|SIEMENS CM VA0  LAB|16|LT|1|CPUIdentificationLabel
0009|SIEMENS CM VA0  LAB|20|LT|1|HeaderVersion
0029|SIEMENS CSA NON-IMAGE|10|OB|1|CSADataInfo
7FE1|SIEMENS CSA NON-IMAGE|10|OB|1|CSAData
0019|SIEMENS CT VA0  COAD|10|DS|1|DistanceSourceToSourceSideCollimator
0019|SIEMENS CT VA0  COAD|11|DS|1|DistanceSourceToDetectorSideCollimator
0019|SIEMENS CT VA0  COAD|20|IS|1|NumberOfPossibleChannels
0019|SIEMENS CT VA0  COAD|21|IS|1|MeanChannelNumber
0019|SIEMENS CT VA0  COAD|22|DS|1|DetectorSpacing
0019|SIEMENS CT VA0  COAD|23|DS|1|DetectorCenter
0019|SIEMENS CT VA0  COAD|24|DS|1|ReadingIntegrationTime
0019|SIEMENS CT VA0  COAD|50|DS|1|DetectorAlignment
0019|SIEMENS CT VA0  COAD|52|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|54|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|60|DS|1|FocusAlignment
0019|SIEMENS CT VA0  COAD|65|UL|1|FocalSpotDeflectionAmplitude
0019|SIEMENS CT VA0  COAD|66|UL|1|FocalSpotDeflectionPhase
0019|SIEMENS CT VA0  COAD|67|UL|1|FocalSpotDeflectionOffset
0019|SIEMENS CT VA0  COAD|70|DS|1|WaterScalingFactor
0019|SIEMENS CT VA0  COAD|71|DS|1|InterpolationFactor
0019|SIEMENS CT VA0  COAD|80|LT|1|PatientRegion
0019|SIEMENS CT VA0  COAD|82|LT|1|PatientPhaseOfLife
0119|MRSC|1181|IS|1|fmSQFitNumber
0019|SIEMENS CT VA0  COAD|94|DS|1|OsteoStandardizationCode
0019|SIEMENS CT VA0  COAD|A3|US|1-n|Unknown
0019|SIEMENS CT VA0  COAD|A4|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|A5|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|A6|US|1-n|Unknown
0019|SIEMENS CT VA0  COAD|A7|US|1-n|Unknown
0019|SIEMENS CT VA0  COAD|A8|US|1-n|Unknown
0019|SIEMENS CT VA0  COAD|A9|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|AA|LT|1|Unknown
0019|SIEMENS CT VA0  COAD|AB|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|AC|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|AD|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|AE|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|AF|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|92|DS|1|OsteoRegressionLineSlope
0019|SIEMENS CT VA0  COAD|93|DS|1|OsteoRegressionLineIntercept
0019|SIEMENS CT VA0  COAD|96|IS|1|OsteoPhantomNumber
0029|SIEMENS CSA HEADER|08|CS|1|CSAImageHeaderType
0029|SIEMENS CSA HEADER|09|LO|1|CSAImageHeaderVersion
0029|SIEMENS CSA HEADER|10|OB|1|CSAImageHeaderInfo
0029|SIEMENS CSA HEADER|18|CS|1|CSASeriesHeaderType
0029|SIEMENS CSA HEADER|19|LO|1|CSASeriesHeaderVersion
0029|SIEMENS CSA HEADER|20|OB|1|CSASeriesHeaderInfo
0029|SIEMENS CSA NON-IMAGE|08|CS|1|CSADataType
0029|SIEMENS CSA NON-IMAGE|09|LO|1|CSADataVersion
0019|SIEMENS CT VA0  COAD|B0|DS|1|FeedPerRotation
0019|SIEMENS CT VA0  COAD|BD|IS|1|PulmoTriggerLevel
0019|SIEMENS CT VA0  COAD|BE|DS|1|ExpiratoricReserveVolume
0019|SIEMENS CT VA0  COAD|BF|DS|1|VitalCapacity
0019|SIEMENS CT VA0  COAD|C0|DS|1|PulmoWater
0019|SIEMENS CT VA0  COAD|C1|DS|1|PulmoAir
0019|SIEMENS CT VA0  COAD|C2|DA|1|PulmoDate
0019|SIEMENS CT VA0  COAD|C3|TM|1|PulmoTime
0019|SIEMENS CT VA0  GEN|10|DS|1|SourceSideCollimatorAperture
0019|SIEMENS CT VA0  GEN|11|DS|1|DetectorSideCollimatorAperture
0019|SIEMENS CT VA0  GEN|20|DS|1|ExposureTime
0019|SIEMENS CT VA0  GEN|21|DS|1|ExposureCurrent
0019|SIEMENS CT VA0  GEN|25|DS|1|KVPGeneratorPowerCurrent
0019|SIEMENS CT VA0  GEN|26|DS|1|GeneratorVoltage
0019|SIEMENS CT VA0  GEN|40|UL|1|MasterControlMask
0019|SIEMENS CT VA0  GEN|42|US|5|ProcessingMask
0019|SIEMENS CT VA0  GEN|44|US|1-n|Unknown
0019|SIEMENS CT VA0  GEN|45|US|1-n|Unknown
0019|SIEMENS CT VA0  GEN|62|IS|1|NumberOfVirtuellChannels
0019|SIEMENS CT VA0  GEN|70|IS|1|NumberOfReadings
0019|SIEMENS CT VA0  GEN|71|LT|1-n|Unknown
0019|SIEMENS CT VA0  GEN|74|IS|1|NumberOfProjections
0019|SIEMENS CT VA0  GEN|75|IS|1|NumberOfBytes
0019|SIEMENS CT VA0  GEN|80|LT|1|ReconstructionAlgorithmSet
0019|SIEMENS CT VA0  GEN|81|LT|1|ReconstructionAlgorithmIndex
0019|SIEMENS CT VA0  GEN|82|LT|1|RegenerationSoftwareVersion
0019|SIEMENS CT VA0  GEN|88|DS|1|Unknown
0021|SIEMENS CT VA0  GEN|10|IS|1|RotationAngle
0021|SIEMENS CT VA0  GEN|11|IS|1|StartAngle
0021|SIEMENS CT VA0  GEN|20|US|1-n|Unknown
0021|SIEMENS CT VA0  GEN|30|IS|1|TopogramTubePosition
0021|SIEMENS CT VA0  GEN|32|DS|1|LengthOfTopogram
0021|SIEMENS CT VA0  GEN|34|DS|1|TopogramCorrectionFactor
0021|SIEMENS CT VA0  GEN|36|DS|1|MaximumTablePosition
0021|SIEMENS CT VA0  GEN|40|IS|1|TableMoveDirectionCode
0021|SIEMENS CT VA0  GEN|45|IS|1|VOIStartRow
0021|SIEMENS CT VA0  GEN|46|IS|1|VOIStopRow
0021|SIEMENS CT VA0  GEN|47|IS|1|VOIStartColumn
0021|SIEMENS CT VA0  GEN|48|IS|1|VOIStopColumn
0021|SIEMENS CT VA0  GEN|49|IS|1|VOIStartSlice
0021|SIEMENS CT VA0  GEN|4a|IS|1|VOIStopSlice
0021|SIEMENS CT VA0  GEN|50|IS|1|VectorStartRow
0021|SIEMENS CT VA0  GEN|51|IS|1|VectorRowStep
0021|SIEMENS CT VA0  GEN|52|IS|1|VectorStartColumn
0021|SIEMENS CT VA0  GEN|53|IS|1|VectorColumnStep
0021|SIEMENS CT VA0  GEN|60|IS|1|RangeTypeCode
0021|SIEMENS CT VA0  GEN|62|IS|1|ReferenceTypeCode
0021|SIEMENS CT VA0  GEN|70|DS|3|ObjectOrientation
0021|SIEMENS CT VA0  GEN|72|DS|3|LightOrientation
0021|SIEMENS CT VA0  GEN|75|DS|1|LightBrightness
0021|SIEMENS CT VA0  GEN|76|DS|1|LightContrast
0021|SIEMENS CT VA0  GEN|7a|IS|2|OverlayThreshold
0021|SIEMENS CT VA0  GEN|7b|IS|2|SurfaceThreshold
0021|SIEMENS CT VA0  GEN|7c|IS|2|GreyScaleThreshold
0021|SIEMENS CT VA0  GEN|a0|DS|1|Unknown
0021|SIEMENS CT VA0  GEN|a2|LT|1|Unknown
0021|SIEMENS CT VA0  GEN|a7|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|10|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|30|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|31|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|32|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|34|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|40|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|42|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|50|LT|1|Unknown
0009|SIEMENS CT VA0  IDE|51|LT|1|Unknown
0009|SIEMENS CT VA0  ORI|20|LT|1|Unknown
0009|SIEMENS CT VA0  ORI|30|LT|1|Unknown
6021|SIEMENS CT VA0  OST|00|LT|1|OsteoContourComment
6021|SIEMENS CT VA0  OST|10|US|256|OsteoContourBuffer
0021|SIEMENS CT VA0  RAW|10|UL|2|CreationMask
0021|SIEMENS CT VA0  RAW|20|UL|2|EvaluationMask
0021|SIEMENS CT VA0  RAW|30|US|7|ExtendedProcessingMask
0021|SIEMENS CT VA0  RAW|40|US|1-n|Unknown
0021|SIEMENS CT VA0  RAW|41|US|1-n|Unknown
0021|SIEMENS CT VA0  RAW|42|US|1-n|Unknown
0021|SIEMENS CT VA0  RAW|43|US|1-n|Unknown
0021|SIEMENS CT VA0  RAW|44|US|1-n|Unknown
0021|SIEMENS CT VA0  RAW|50|LT|1|Unknown
0009|SIEMENS DICOM|10|UN|1|Unknown
0009|SIEMENS DICOM|12|LT|1|Unknown
0019|SIEMENS DLR.01|10|LT|1|MeasurementMode
0019|SIEMENS DLR.01|11|LT|1|ImageType
0019|SIEMENS DLR.01|15|LT|1|SoftwareVersion
0019|SIEMENS DLR.01|20|LT|1|MPMCode
0019|SIEMENS DLR.01|21|LT|1|Latitude
0019|SIEMENS DLR.01|22|LT|1|Sensitivity
0019|SIEMENS DLR.01|23|LT|1|EDR
0019|SIEMENS DLR.01|24|LT|1|LFix
0019|SIEMENS DLR.01|25|LT|1|SFix
0019|SIEMENS DLR.01|26|LT|1|PresetMode
0019|SIEMENS DLR.01|27|LT|1|Region
0019|SIEMENS DLR.01|28|LT|1|Subregion
0019|SIEMENS DLR.01|30|LT|1|Orientation
0019|SIEMENS DLR.01|31|LT|1|MarkOnFilm
0019|SIEMENS DLR.01|32|LT|1|RotationOnDRC
0019|SIEMENS DLR.01|40|LT|1|ReaderType
0019|SIEMENS DLR.01|41|LT|1|SubModality
0019|SIEMENS DLR.01|42|LT|1|ReaderSerialNumber
0019|SIEMENS DLR.01|50|LT|1|CassetteScale
0019|SIEMENS DLR.01|51|LT|1|CassetteMatrix
0019|SIEMENS DLR.01|52|LT|1|CassetteSubmatrix
0019|SIEMENS DLR.01|53|LT|1|Barcode
0019|SIEMENS DLR.01|60|LT|1|ContrastType
0019|SIEMENS DLR.01|61|LT|1|RotationAmount
0019|SIEMENS DLR.01|62|LT|1|RotationCenter
0019|SIEMENS DLR.01|63|LT|1|DensityShift
0019|SIEMENS DLR.01|64|US|1|FrequencyRank
0019|SIEMENS DLR.01|65|LT|1|FrequencyEnhancement
0019|SIEMENS DLR.01|66|LT|1|FrequencyType
0019|SIEMENS DLR.01|67|LT|1|KernelLength
0019|SIEMENS DLR.01|68|UL|1|KernelMode
0019|SIEMENS DLR.01|69|UL|1|ConvolutionMode
0019|SIEMENS DLR.01|70|LT|1|PLASource
0019|SIEMENS DLR.01|71|LT|1|PLADestination
0019|SIEMENS DLR.01|75|LT|1|UIDOriginalImage
0019|SIEMENS DLR.01|76|LT|1|Unknown
0019|SIEMENS DLR.01|80|LT|1|ReaderHeader
0019|SIEMENS DLR.01|90|LT|1|PLAOfSecondaryDestination
0019|SIEMENS DLR.01|a0|DS|1|Unknown
0019|SIEMENS DLR.01|a1|DS|1|Unknown
0041|SIEMENS DLR.01|10|US|1|NumberOfHardcopies
0041|SIEMENS DLR.01|20|LT|1|FilmFormat
0041|SIEMENS DLR.01|30|LT|1|FilmSize
0041|SIEMENS DLR.01|31|LT|1|FullFilmFormat
0003|SIEMENS ISI|08|US|1|ISICommandField
0003|SIEMENS ISI|11|US|1|AttachIDApplicationCode
0003|SIEMENS ISI|12|UL|1|AttachIDMessageCount
0003|SIEMENS ISI|13|DA|1|AttachIDDate
0003|SIEMENS ISI|14|TM|1|AttachIDTime
0003|SIEMENS ISI|20|US|1|MessageType
0003|SIEMENS ISI|30|DA|1|MaxWaitingDate
0003|SIEMENS ISI|31|TM|1|MaxWaitingTime
0009|SIEMENS ISI|01|UN|1|RISPatientInfoIMGEF
0011|SIEMENS ISI|03|LT|1|PatientUID
0011|SIEMENS ISI|04|LT|1|PatientID
0011|SIEMENS ISI|0a|LT|1|CaseID
0011|SIEMENS ISI|22|LT|1|RequestID
0011|SIEMENS ISI|23|LT|1|ExaminationUID
0011|SIEMENS ISI|a1|DA|1|PatientRegistrationDate
0011|SIEMENS ISI|a2|TM|1|PatientRegistrationTime
0011|SIEMENS ISI|b0|LT|1|PatientLastName
0011|SIEMENS ISI|b2|LT|1|PatientFirstName
0011|SIEMENS ISI|b4|LT|1|PatientHospitalStatus
0011|SIEMENS ISI|bc|TM|1|CurrentLocationTime
0011|SIEMENS ISI|c0|LT|1|PatientInsuranceStatus
0011|SIEMENS ISI|d0|LT|1|PatientBillingType
0011|SIEMENS ISI|d2|LT|1|PatientBillingAddress
0031|SIEMENS ISI|12|LT|1|ExaminationReason
0031|SIEMENS ISI|30|DA|1|RequestedDate
0031|SIEMENS ISI|32|TM|1|WorklistRequestStartTime
0031|SIEMENS ISI|33|TM|1|WorklistRequestEndTime
0031|SIEMENS ISI|4a|TM|1|RequestedTime
0031|SIEMENS ISI|80|LT|1|RequestedLocation
0055|SIEMENS ISI|46|LT|1|CurrentWard
0193|SIEMENS ISI|02|DS|1|RISKey
0307|SIEMENS ISI|01|UN|1|RISWorklistIMGEF
0309|SIEMENS ISI|01|UN|1|RISReportIMGEF
4009|SIEMENS ISI|01|LT|1|ReportID
4009|SIEMENS ISI|20|LT|1|ReportStatus
4009|SIEMENS ISI|30|DA|1|ReportCreationDate
4009|SIEMENS ISI|70|LT|1|ReportApprovingPhysician
4009|SIEMENS ISI|e0|LT|1|ReportText
4009|SIEMENS ISI|e1|LT|1|ReportAuthor
4009|SIEMENS ISI|e3|LT|1|ReportingRadiologist
0029|SIEMENS MED DISPLAY|04|LT|1|PhotometricInterpretation
0029|SIEMENS MED DISPLAY|10|US|1|RowsOfSubmatrix
0029|SIEMENS MED DISPLAY|11|US|1|ColumnsOfSubmatrix
0029|SIEMENS MED DISPLAY|20|US|1|Unknown
0029|SIEMENS MED DISPLAY|21|US|1|Unknown
0029|SIEMENS MED DISPLAY|50|US|1|OriginOfSubmatrix
0029|SIEMENS MED DISPLAY|99|LT|1|ShutterType
0029|SIEMENS MED DISPLAY|a0|US|1|RowsOfRectangularShutter
0029|SIEMENS MED DISPLAY|a1|US|1|ColumnsOfRectangularShutter
0029|SIEMENS MED DISPLAY|a2|US|1|OriginOfRectangularShutter
0029|SIEMENS MED DISPLAY|b0|US|1|RadiusOfCircularShutter
0029|SIEMENS MED DISPLAY|b2|US|1|OriginOfCircularShutter
0029|SIEMENS MED DISPLAY|c1|US|1|ContourOfIrregularShutter
0029|SIEMENS MED HG|10|US|1|ListOfGroupNumbers
0029|SIEMENS MED HG|15|LT|1|ListOfShadowOwnerCodes
0029|SIEMENS MED HG|20|US|1|ListOfElementNumbers
0029|SIEMENS MED HG|30|US|1|ListOfTotalDisplayLength
0029|SIEMENS MED HG|40|LT|1|ListOfDisplayPrefix
0029|SIEMENS MED HG|50|LT|1|ListOfDisplayPostfix
0029|SIEMENS MED HG|60|US|1|ListOfTextPosition
0029|SIEMENS MED HG|70|LT|1|ListOfTextConcatenation
0029|SIEMENS MED MG|10|US|1|ListOfGroupNumbers
0029|SIEMENS MED MG|15|LT|1|ListOfShadowOwnerCodes
0029|SIEMENS MED MG|20|US|1|ListOfElementNumbers
0029|SIEMENS MED MG|30|US|1|ListOfTotalDisplayLength
0029|SIEMENS MED MG|40|LT|1|ListOfDisplayPrefix
0029|SIEMENS MED MG|50|LT|1|ListOfDisplayPostfix
0029|SIEMENS MED MG|60|US|1|ListOfTextPosition
0029|SIEMENS MED MG|70|LT|1|ListOfTextConcatenation
0009|SIEMENS MED|10|LO|1|RecognitionCode
0009|SIEMENS MED|30|UL|1|ByteOffsetOfOriginalHeader
0009|SIEMENS MED|31|UL|1|LengthOfOriginalHeader
0009|SIEMENS MED|40|UL|1|ByteOffsetOfPixelmatrix
0009|SIEMENS MED|41|UL|1|LengthOfPixelmatrixInBytes
0009|SIEMENS MED|50|LT|1|Unknown
0009|SIEMENS MED|51|LT|1|Unknown
0009|SIEMENS MED|f5|LT|1|PDMEFIDPlaceholder
0009|SIEMENS MED|f6|LT|1|PDMDataObjectTypeExtension
0021|SIEMENS MED|10|DS|1|Zoom
0021|SIEMENS MED|12|IS|1|TubeAngle
0021|SIEMENS MED|20|US|1|ROIMask
7001|SIEMENS MED|10|LT|1|Dummy
7003|SIEMENS MED|10|LT|1|Header
7005|SIEMENS MED|10|LT|1|Dummy
0119|MRSC|11a0|CS|1|PhantCalibType
0029|SIEMENS MEDCOM HEADER|09|LO|1|MedComHeaderVersion
0029|SIEMENS MEDCOM HEADER|10|OB|1|MedComHeaderInfo
0029|SIEMENS MEDCOM HEADER|20|OB|1|MedComHistoryInformation
0029|SIEMENS MEDCOM HEADER|31|LO|1|PMTFInformation1
0029|SIEMENS MEDCOM HEADER|32|UL|1|PMTFInformation2
0029|SIEMENS MEDCOM HEADER|33|UL|1|PMTFInformation3
0029|SIEMENS MEDCOM HEADER|34|CS|1|PMTFInformation4
0029|SIEMENS MEDCOM HEADER|35|UL|1|PMTFInformation5
0029|SIEMENS MEDCOM HEADER|40|SQ|1|ApplicationHeaderSequence
0029|SIEMENS MEDCOM HEADER|41|CS|1|ApplicationHeaderType
0029|SIEMENS MEDCOM HEADER|42|LO|1|ApplicationHeaderID
0019|SIEMENS MR VA0  COAD|12|DS|1|MagneticFieldStrength
0019|SIEMENS MR VA0  COAD|14|DS|1|ADCVoltage
0019|SIEMENS MR VA0  COAD|16|DS|2|ADCOffset
0019|SIEMENS MR VA0  COAD|20|DS|1|TransmitterAmplitude
0019|SIEMENS MR VA0  COAD|21|IS|1|NumberOfTransmitterAmplitudes
0019|SIEMENS MR VA0  COAD|22|DS|1|TransmitterAttenuator
0019|SIEMENS MR VA0  COAD|24|DS|1|TransmitterCalibration
0019|SIEMENS MR VA0  COAD|26|DS|1|TransmitterReference
0019|SIEMENS MR VA0  COAD|50|DS|1|ReceiverTotalGain
0019|SIEMENS MR VA0  COAD|51|DS|1|ReceiverAmplifierGain
0019|SIEMENS MR VA0  COAD|52|DS|1|ReceiverPreamplifierGain
0019|SIEMENS MR VA0  COAD|54|DS|1|ReceiverCableAttenuation
0019|SIEMENS MR VA0  COAD|55|DS|1|ReceiverReferenceGain
0019|SIEMENS MR VA0  COAD|56|DS|1|ReceiverFilterFrequency
0019|SIEMENS MR VA0  COAD|60|DS|1|ReconstructionScaleFactor
0019|SIEMENS MR VA0  COAD|62|DS|1|ReferenceScaleFactor
0019|SIEMENS MR VA0  COAD|70|DS|1|PhaseGradientAmplitude
0019|SIEMENS MR VA0  COAD|71|DS|1|ReadoutGradientAmplitude
0019|SIEMENS MR VA0  COAD|72|DS|1|SelectionGradientAmplitude
0019|SIEMENS MR VA0  COAD|80|DS|3|GradientDelayTime
0019|SIEMENS MR VA0  COAD|82|DS|1|TotalGradientDelayTime
0019|SIEMENS MR VA0  COAD|90|LT|1|SensitivityCorrectionLabel
0019|SIEMENS MR VA0  COAD|91|DS|6|SaturationPhaseEncodingVectorCoronalComponent
0019|SIEMENS MR VA0  COAD|92|DS|6|SaturationReadoutVectorCoronalComponent
0019|SIEMENS MR VA0  COAD|a0|US|3|RFWatchdogMask
0019|SIEMENS MR VA0  COAD|a1|DS|1|EPIReconstructionSlope
0019|SIEMENS MR VA0  COAD|a2|DS|1|RFPowerErrorIndicator
0019|SIEMENS MR VA0  COAD|a5|DS|3|SpecificAbsorptionRateWholeBody
0019|SIEMENS MR VA0  COAD|a6|DS|3|SpecificEnergyDose
0019|SIEMENS MR VA0  COAD|b0|UL|1|AdjustmentStatusMask
0019|SIEMENS MR VA0  COAD|c1|DS|6|EPICapacity
0019|SIEMENS MR VA0  COAD|c2|DS|3|EPIInductance
0019|SIEMENS MR VA0  COAD|c3|IS|1-n|EPISwitchConfigurationCode
0019|SIEMENS MR VA0  COAD|c4|IS|1-n|EPISwitchHardwareCode
0019|SIEMENS MR VA0  COAD|c5|DS|1-n|EPISwitchDelayTime
0019|SIEMENS MR VA0  COAD|d1|DS|1|FlowSensitivity
0019|SIEMENS MR VA0  COAD|d2|LT|1|CalculationSubmode
0029|SIEMENS MEDCOM HEADER|44|OB|1|ApplicationHeaderInfo
0029|SIEMENS MEDCOM HEADER|50|LO|8|WorkflowControlFlags
0029|SIEMENS MEDCOM HEADER|51|CS|1|ArchiveManagementFlagKeepOnline
0029|SIEMENS MEDCOM HEADER|52|CS|1|ArchiveManagementFlagDoNotArchive
0029|SIEMENS MEDCOM HEADER|53|CS|1|ImageLocationStatus
0029|SIEMENS MEDCOM HEADER|54|DS|1|EstimatedRetrieveTime
0029|SIEMENS MEDCOM HEADER|55|DS|1|DataSizeOfRetrievedImages
0029|SIEMENS MEDCOM HEADER2|60|LO|1|SeriesWorkflowStatus
0029|SIEMENS MEDCOM OOG|08|CS|1|MEDCOMOOGType
0029|SIEMENS MEDCOM OOG|09|LO|1|MEDCOMOOGVersion
0029|SIEMENS MEDCOM OOG|10|OB|1|MEDCOMOOGInfo
0019|SIEMENS MR VA0  COAD|d3|DS|1|FieldOfViewRatio
0019|SIEMENS MR VA0  COAD|d4|IS|1|BaseRawMatrixSize
0019|SIEMENS MR VA0  COAD|d5|IS|1|2DOversamplingLines
0019|SIEMENS MR VA0  COAD|d6|IS|1|3DPhaseOversamplingPartitions
0019|SIEMENS MR VA0  COAD|d7|IS|1|EchoLinePosition
0019|SIEMENS MR VA0  COAD|d8|IS|1|EchoColumnPosition
0019|SIEMENS MR VA0  COAD|d9|IS|1|LinesPerSegment
0019|SIEMENS MR VA0  COAD|da|LT|1|PhaseCodingDirection
0019|SIEMENS MR VA0  GEN|10|DS|1|TotalMeasurementTimeNominal
0019|SIEMENS MR VA0  GEN|11|DS|1|TotalMeasurementTimeCurrent
0019|SIEMENS MR VA0  GEN|12|DS|1|StartDelayTime
0019|SIEMENS MR VA0  GEN|13|DS|1|DwellTime
0019|SIEMENS MR VA0  GEN|14|IS|1|NumberOfPhases
0019|SIEMENS MR VA0  GEN|16|UL|2|SequenceControlMask
0019|SIEMENS MR VA0  GEN|18|UL|1|MeasurementStatusMask
0019|SIEMENS MR VA0  GEN|20|IS|1|NumberOfFourierLinesNominal
0019|SIEMENS MR VA0  GEN|21|IS|1|NumberOfFourierLinesCurrent
0019|SIEMENS MR VA0  GEN|26|IS|1|NumberOfFourierLinesAfterZero
0019|SIEMENS MR VA0  GEN|28|IS|1|FirstMeasuredFourierLine
0019|SIEMENS MR VA0  GEN|30|IS|1|AcquisitionColumns
0019|SIEMENS MR VA0  GEN|31|IS|1|ReconstructionColumns
0019|SIEMENS MR VA0  GEN|40|IS|1|ArrayCoilElementNumber
0019|SIEMENS MR VA0  GEN|41|UL|1|ArrayCoilElementSelectMask
0019|SIEMENS MR VA0  GEN|42|UL|1|ArrayCoilElementDataMask
0019|SIEMENS MR VA0  GEN|43|IS|1-n|ArrayCoilElementToADCConnect
0019|SIEMENS MR VA0  GEN|44|DS|1-n|ArrayCoilElementNoiseLevel
0019|SIEMENS MR VA0  GEN|45|IS|1|ArrayCoilADCPairNumber
0019|SIEMENS MR VA0  GEN|46|UL|1|ArrayCoilCombinationMask
0019|SIEMENS MR VA0  GEN|50|IS|1|NumberOfAverages
0019|SIEMENS MR VA0  GEN|60|DS|1|FlipAngle
0019|SIEMENS MR VA0  GEN|70|IS|1|NumberOfPrescans
0019|SIEMENS MR VA0  GEN|81|LT|1|FilterTypeForRawData
0019|SIEMENS MR VA0  GEN|82|DS|1-n|FilterParameterForRawData
0019|SIEMENS MR VA0  GEN|83|LT|1|FilterTypeForImageData
0019|SIEMENS MR VA0  GEN|84|DS|1-n|FilterParameterForImageData
0019|SIEMENS MR VA0  GEN|85|LT|1|FilterTypeForPhaseCorrection
0019|SIEMENS MR VA0  GEN|86|DS|1-n|FilterParameterForPhaseCorrection
0019|SIEMENS MR VA0  GEN|87|LT|1|NormalizationFilterTypeForImageData
0019|SIEMENS MR VA0  GEN|88|DS|1-n|NormalizationFilterParameterForImageData
0019|SIEMENS MR VA0  GEN|90|IS|1|NumberOfSaturationRegions
0019|SIEMENS MR VA0  GEN|91|DS|6|SaturationPhaseEncodingVectorSagittalComponent
0019|SIEMENS MR VA0  GEN|92|DS|6|SaturationReadoutVectorSagittalComponent
0019|SIEMENS MR VA0  GEN|93|DS|1|EPIStimulationMonitorMode
0019|SIEMENS MR VA0  GEN|94|DS|1|ImageRotationAngle
0019|SIEMENS MR VA0  GEN|96|UL|3|CoilIDMask
0019|SIEMENS MR VA0  GEN|97|UL|2|CoilClassMask
0019|SIEMENS MR VA0  GEN|98|DS|3|CoilPosition
0019|SIEMENS MR VA0  GEN|a0|DS|1|EPIReconstructionPhase
0019|SIEMENS MR VA0  GEN|a1|DS|1|EPIReconstructionSlope
0021|SIEMENS MR VA0  GEN|20|IS|1|PhaseCorrectionRowsSequence
0021|SIEMENS MR VA0  GEN|21|IS|1|PhaseCorrectionColumnsSequence
0021|SIEMENS MR VA0  GEN|22|IS|1|PhaseCorrectionRowsReconstruction
0021|SIEMENS MR VA0  GEN|24|IS|1|PhaseCorrectionColumnsReconstruction
0021|SIEMENS MR VA0  GEN|30|IS|1|NumberOf3DRawPartitionsNominal
0021|SIEMENS MR VA0  GEN|31|IS|1|NumberOf3DRawPartitionsCurrent
0021|SIEMENS MR VA0  GEN|34|IS|1|NumberOf3DImagePartitions
0021|SIEMENS MR VA0  GEN|36|IS|1|Actual3DImagePartitionNumber
0021|SIEMENS MR VA0  GEN|39|DS|1|SlabThickness
0021|SIEMENS MR VA0  GEN|40|IS|1|NumberOfSlicesNominal
0021|SIEMENS MR VA0  GEN|41|IS|1|NumberOfSlicesCurrent
0021|SIEMENS MR VA0  GEN|42|IS|1|CurrentSliceNumber
0021|SIEMENS MR VA0  GEN|43|IS|1|CurrentGroupNumber
0021|SIEMENS MR VA0  GEN|44|DS|1|CurrentSliceDistanceFactor
0021|SIEMENS MR VA0  GEN|45|IS|1|MIPStartRow
0021|SIEMENS MR VA0  GEN|46|IS|1|MIPStopRow
0021|SIEMENS MR VA0  GEN|47|IS|1|MIPStartColumn
0021|SIEMENS MR VA0  GEN|48|IS|1|MIPStartColumn
0021|SIEMENS MR VA0  GEN|49|IS|1|MIPStartSlice Name=
0021|SIEMENS MR VA0  GEN|4a|IS|1|MIPStartSlice
0021|SIEMENS MR VA0  GEN|4f|LT|1|OrderofSlices
0021|SIEMENS MR VA0  GEN|50|US|1|SignalMask
0021|SIEMENS MR VA0  GEN|52|DS|1|DelayAfterTrigger
0021|SIEMENS MR VA0  GEN|53|IS|1|RRInterval
0021|SIEMENS MR VA0  GEN|54|DS|1|NumberOfTriggerPulses
0021|SIEMENS MR VA0  GEN|56|DS|1|RepetitionTimeEffective
0021|SIEMENS MR VA0  GEN|57|LT|1|GatePhase
0021|SIEMENS MR VA0  GEN|58|DS|1|GateThreshold
0021|SIEMENS MR VA0  GEN|59|DS|1|GatedRatio
0021|SIEMENS MR VA0  GEN|60|IS|1|NumberOfInterpolatedImages
0021|SIEMENS MR VA0  GEN|70|IS|1|NumberOfEchoes
0021|SIEMENS MR VA0  GEN|72|DS|1|SecondEchoTime
0021|SIEMENS MR VA0  GEN|73|DS|1|SecondRepetitionTime
0021|SIEMENS MR VA0  GEN|80|IS|1|CardiacCode
0021|SIEMENS MR VA0  GEN|91|DS|6|SaturationPhaseEncodingVectorTransverseComponent
0021|SIEMENS MR VA0  GEN|92|DS|6|SaturationReadoutVectorTransverseComponent
0021|SIEMENS MR VA0  GEN|93|DS|1|EPIChangeValueOfMagnitude
0021|SIEMENS MR VA0  GEN|94|DS|1|EPIChangeValueOfXComponent
0021|SIEMENS MR VA0  GEN|95|DS|1|EPIChangeValueOfYComponent
0021|SIEMENS MR VA0  GEN|96|DS|1|EPIChangeValueOfZComponent
0021|SIEMENS MR VA0  RAW|00|LT|1|SequenceType
0021|SIEMENS MR VA0  RAW|01|IS|1|VectorSizeOriginal
0021|SIEMENS MR VA0  RAW|02|IS|1|VectorSizeExtended
0021|SIEMENS MR VA0  RAW|03|DS|1|AcquiredSpectralRange
0021|SIEMENS MR VA0  RAW|04|DS|3|VOIPosition
0021|SIEMENS MR VA0  RAW|05|DS|3|VOISize
0021|SIEMENS MR VA0  RAW|06|IS|3|CSIMatrixSizeOriginal
0021|SIEMENS MR VA0  RAW|07|IS|3|CSIMatrixSizeExtended
0021|SIEMENS MR VA0  RAW|08|DS|3|SpatialGridShift
0021|SIEMENS MR VA0  RAW|09|DS|1|SignalLimitsMinimum
0019|SVISION|81|IS|1|ObjectPosition
0021|SIEMENS MR VA0  RAW|10|DS|1|SignalLimitsMaximum
0021|SIEMENS MR VA0  RAW|11|DS|1|SpecInfoMask
0021|SIEMENS MR VA0  RAW|12|DS|1|EPITimeRateOfChangeOfMagnitude
0021|SIEMENS MR VA0  RAW|13|DS|1|EPITimeRateOfChangeOfXComponent
0021|SIEMENS MR VA0  RAW|14|DS|1|EPITimeRateOfChangeOfYComponent
0021|SIEMENS MR VA0  RAW|15|DS|1|EPITimeRateOfChangeOfZComponent
0021|SIEMENS MR VA0  RAW|16|DS|1|EPITimeRateOfChangeLegalLimit1
0021|SIEMENS MR VA0  RAW|17|DS|1|EPIOperationModeFlag
0021|SIEMENS MR VA0  RAW|18|DS|1|EPIFieldCalculationSafetyFactor
0021|SIEMENS MR VA0  RAW|19|DS|1|EPILegalLimit1OfChangeValue
0021|SIEMENS MR VA0  RAW|20|DS|1|EPILegalLimit2OfChangeValue
0021|SIEMENS MR VA0  RAW|21|DS|1|EPIRiseTime
0021|SIEMENS MR VA0  RAW|30|DS|16|ArrayCoilADCOffset
0021|SIEMENS MR VA0  RAW|31|DS|16|ArrayCoilPreamplifierGain
0021|SIEMENS MR VA0  RAW|50|LT|1|SaturationType
0021|SIEMENS MR VA0  RAW|51|DS|3|SaturationNormalVector
0021|SIEMENS MR VA0  RAW|52|DS|3|SaturationPositionVector
0021|SIEMENS MR VA0  RAW|53|DS|6|SaturationThickness
0021|SIEMENS MR VA0  RAW|54|DS|6|SaturationWidth
0021|SIEMENS MR VA0  RAW|55|DS|6|SaturationDistance
7fe3|SIEMENS NUMARIS II|00|LT|1|ImageGraphicsFormatCode
7fe3|SIEMENS NUMARIS II|10|OB|1|ImageGraphics
7fe3|SIEMENS NUMARIS II|20|OB|1|ImageGraphicsDummy
0011|SIEMENS RA GEN|20|SL|1|FluoroTimer
0011|SIEMENS RA GEN|25|SL|1|PtopDoseAreaProduct
0011|SIEMENS RA GEN|26|SL|1|PtopTotalSkinDose
0011|SIEMENS RA GEN|30|LT|1|Unknown
0011|SIEMENS RA GEN|35|LO|1|PatientInitialPuckCounter
0011|SIEMENS RA GEN|40|SS|1|SPIDataObjectType
0019|SIEMENS RA GEN|15|LO|1|AcquiredPlane
0019|SIEMENS RA GEN|1f|SS|1|DefaultTableIsoCenterHeight
0019|SIEMENS RA GEN|20|SL|1|SceneFlag
0019|SIEMENS RA GEN|22|SL|1|RefPhotofileFlag
0019|SIEMENS RA GEN|24|LO|1|SceneName
0019|SIEMENS RA GEN|26|SS|1|AcquisitionIndex
0019|SIEMENS RA GEN|28|SS|1|MixedPulseMode
0019|SIEMENS RA GEN|2a|SS|1|NoOfPositions
0019|SIEMENS RA GEN|2c|SS|1|NoOfPhases
0019|SIEMENS RA GEN|2e|SS|1-n|FrameRateForPositions
0019|SIEMENS RA GEN|30|SS|1-n|NoOfFramesForPositions
0019|SIEMENS RA GEN|32|SS|1|SteppingDirection
0019|SIEMENS RA GEN|34|US|1|Unknown
0019|SIEMENS RA GEN|36|US|1|Unknown
0019|SIEMENS RA GEN|38|US|1|Unknown
0019|SIEMENS RA GEN|3a|US|1|Unknown
0019|SIEMENS RA GEN|3c|US|1|Unknown
0019|SIEMENS RA GEN|3e|US|1|Unknown
0019|SIEMENS RA GEN|40|US|1|Unknown
0019|SIEMENS RA GEN|42|US|1|Unknown
0019|SIEMENS RA GEN|44|SS|1|ImageTransferDelay
0019|SIEMENS RA GEN|46|SL|1|InversFlag
0019|SIEMENS RA GEN|48|US|1|Unknown
0019|SIEMENS RA GEN|4a|US|1|Unknown
0019|SIEMENS RA GEN|4c|SS|1|BlankingCircleDiameter
0019|SIEMENS RA GEN|50|SL|1|StandDataValid
0019|SIEMENS RA GEN|54|SS|1|TableAxisRotation
0019|SIEMENS RA GEN|56|SS|1|TableLongitudalPosition
0019|SIEMENS RA GEN|58|SS|1|TableSideOffset
0019|SIEMENS RA GEN|5a|SS|1|TableIsoCenterHeight
0019|SIEMENS RA GEN|5c|UN|1|Unknown
0019|SIEMENS RA GEN|5e|SL|1|CollimationDataValid
0019|SIEMENS RA GEN|60|SL|1|PeriSequenceNo
0019|SIEMENS RA GEN|62|SL|1|PeriTotalScenes
0019|SIEMENS RA GEN|64|SL|1|PeriOverlapTop
0019|SIEMENS RA GEN|66|SL|1|PeriOverlapBottom
0019|SIEMENS RA GEN|68|SL|1|RawImageNumber
0019|SIEMENS RA GEN|6a|SL|1|XRayDataValid
0019|SIEMENS RA GEN|70|US|1-n|Unknown
0019|SIEMENS RA GEN|72|US|1-n|Unknown
0019|SIEMENS RA GEN|74|US|1-n|Unknown
0019|SIEMENS RA GEN|76|SL|1|FillingAverageFactor
0019|SIEMENS RA GEN|78|US|1-n|Unknown
0019|SIEMENS RA GEN|7a|US|1-n|Unknown
0019|SIEMENS RA GEN|7c|US|1-n|Unknown
0019|SIEMENS RA GEN|7e|US|1-n|Unknown
0019|SIEMENS RA GEN|80|US|1-n|Unknown
0019|SIEMENS RA GEN|82|US|1-n|Unknown
0019|SIEMENS RA GEN|84|US|1-n|Unknown
0019|SIEMENS RA GEN|86|US|1-n|Unknown
0019|SIEMENS RA GEN|88|US|1-n|Unknown
0019|SIEMENS RA GEN|8a|US|1-n|Unknown
0019|SIEMENS RA GEN|8c|US|1-n|Unknown
0019|SIEMENS RA GEN|8e|US|1-n|Unknown
0019|SIEMENS RA GEN|92|US|1-n|Unknown
0019|SIEMENS RA GEN|94|US|1-n|Unknown
0019|SIEMENS RA GEN|96|US|1-n|Unknown
0019|SIEMENS RA GEN|98|US|1-n|Unknown
0019|SIEMENS RA GEN|9a|US|1-n|Unknown
0019|SIEMENS RA GEN|9c|SL|1|IntensifierLevelCalibrationFactor
0019|SIEMENS RA GEN|9e|SL|1|NativeReviewFlag
0019|SIEMENS RA GEN|a2|SL|1|SceneNumber
0019|SIEMENS RA GEN|a4|SS|1|AcquisitionMode
0019|SIEMENS RA GEN|a5|SS|1|AcquisitonFrameRate
0019|SIEMENS RA GEN|a6|SL|1|ECGFlag
0019|SIEMENS RA GEN|a7|SL|1|AdditionalSceneData
0019|SIEMENS RA GEN|a8|SL|1|FileCopyFlag
0019|SIEMENS RA GEN|a9|SL|1|PhlebovisionFlag
0019|SIEMENS RA GEN|aa|SL|1|Co2Flag
0019|SIEMENS RA GEN|ab|SS|1|MaxSpeed
0019|SIEMENS RA GEN|ac|SS|1|StepWidth
0019|SIEMENS RA GEN|ad|SL|1|DigitalAcquisitionZoom
0019|SIEMENS RA GEN|ff|SS|1-n|Internal
0021|SIEMENS RA GEN|15|SS|1|ImagesInStudy
0021|SIEMENS RA GEN|20|SS|1|ScenesInStudy
0021|SIEMENS RA GEN|25|SS|1|ImagesInPhotofile
0021|SIEMENS RA GEN|27|SS|1|PlaneBImagesExist
0021|SIEMENS RA GEN|28|SS|1|NoOf2MBChunks
0021|SIEMENS RA GEN|30|SS|1|ImagesInAllScenes
0021|SIEMENS RA GEN|40|SS|1|ArchiveSWInternalVersion
0011|SIEMENS RA PLANE A|28|SL|1|FluoroTimerA
0011|SIEMENS RA PLANE A|29|SL|1|FluoroSkinDoseA
0011|SIEMENS RA PLANE A|2a|SL|1|TotalSkinDoseA
0011|SIEMENS RA PLANE A|2b|SL|1|FluoroDoseAreaProductA
0011|SIEMENS RA PLANE A|2c|SL|1|TotalDoseAreaProductA
0019|SIEMENS RA PLANE A|15|LT|1|OfflineUID
0019|SIEMENS RA PLANE A|18|SS|1|Internal
0019|SIEMENS RA PLANE A|19|SS|1|Internal
0019|SIEMENS RA PLANE A|1a|SS|1|Internal
0019|SIEMENS RA PLANE A|1b|SS|1|Internal
0019|SIEMENS RA PLANE A|1c|SS|1|Internal
0019|SIEMENS RA PLANE A|1d|SS|1|Internal
0019|SIEMENS RA PLANE A|1e|SS|1|Internal
0019|SIEMENS RA PLANE A|1f|SS|1-n|Internal
0019|SIEMENS RA PLANE A|20|SS|1|SystemCalibFactorPlaneA
0019|SIEMENS RA PLANE A|22|SS|1|XRayParameterSetNo
0019|SIEMENS RA PLANE A|24|SS|1|XRaySystem
0019|SIEMENS RA PLANE A|26|US|1|Unknown
0019|SIEMENS RA PLANE A|28|SS|1|AcquiredDisplayMode
0019|SIEMENS RA PLANE A|2a|SS|1|AcquisitionDelay
0019|SIEMENS RA PLANE A|2c|US|1|Unknown
0019|SIEMENS RA PLANE A|2e|SS|1|MaxFramesLimit
0019|SIEMENS RA PLANE A|30|US|1|MaximumFrameSizeNIU
0019|SIEMENS RA PLANE A|32|SS|1|SubtractedFilterType
0019|SIEMENS RA PLANE A|34|SS|1|FilterFactorNative
0019|SIEMENS RA PLANE A|36|SS|1|AnatomicBackgroundFactor
0019|SIEMENS RA PLANE A|38|SS|1|WindowUpperLimitNative
0019|SIEMENS RA PLANE A|3a|SS|1|WindowLowerLimitNative
0019|SIEMENS RA PLANE A|3c|SS|1|WindowBrightnessPhase1
0019|SIEMENS RA PLANE A|3e|SS|1|WindowBrightnessPhase2
0019|SIEMENS RA PLANE A|40|SS|1|WindowContrastPhase1
0019|SIEMENS RA PLANE A|42|SS|1|WindowContrastPhase2
0019|SIEMENS RA PLANE A|44|SS|1|FilterFactorSub
0019|SIEMENS RA PLANE A|46|SS|1|PeakOpacified
0019|SIEMENS RA PLANE A|48|SL|1|MaskFrame
0019|SIEMENS RA PLANE A|4a|SL|1|BIHFrame
0019|SIEMENS RA PLANE A|4c|SS|1|CentBeamAngulationCaudCran
0019|SIEMENS RA PLANE A|4e|SS|1|CentBeamAngulationLRAnterior
0019|SIEMENS RA PLANE A|50|SS|1|LongitudinalPosition
0019|SIEMENS RA PLANE A|52|SS|1|SideOffset
0019|SIEMENS RA PLANE A|54|SS|1|IsoCenterHeight
0019|SIEMENS RA PLANE A|56|SS|1|ImageTwist
0019|SIEMENS RA PLANE A|58|SS|1|SourceImageDistance
0019|SIEMENS RA PLANE A|5a|SS|1|MechanicalMagnificationFactor
0019|SIEMENS RA PLANE A|5c|SL|1|CalibrationFlag
0019|SIEMENS RA PLANE A|5e|SL|1|CalibrationAngleCranCaud
0019|SIEMENS RA PLANE A|60|SL|1|CalibrationAngleRAOLAO
0019|SIEMENS RA PLANE A|62|SL|1|CalibrationTableToFloorDist
0019|SIEMENS RA PLANE A|64|SL|1|CalibrationIsocenterToFloorDist
0019|SIEMENS RA PLANE A|66|SL|1|CalibrationIsocenterToSourceDist
0019|SIEMENS RA PLANE A|68|SL|1|CalibrationSourceToII
0019|SIEMENS RA PLANE A|6a|SL|1|CalibrationIIZoom
0019|SIEMENS RA PLANE A|6c|SL|1|CalibrationIIField
0019|SIEMENS RA PLANE A|6e|SL|1|CalibrationFactor
0019|SIEMENS RA PLANE A|70|SL|1|CalibrationObjectToImageDistance
0019|SIEMENS RA PLANE A|72|SL|1-n|CalibrationSystemFactor
0019|SIEMENS RA PLANE A|74|SL|1-n|CalibrationSystemCorrection
0019|SIEMENS RA PLANE A|76|SL|1-n|CalibrationSystemIIFormats
0019|SIEMENS RA PLANE A|78|SL|1|CalibrationGantryDataValid
0019|SIEMENS RA PLANE A|7a|SS|1|CollimatorSquareBreadth
0019|SIEMENS RA PLANE A|7c|SS|1|CollimatorSquareHeight
0019|SIEMENS RA PLANE A|7e|SS|1|CollimatorSquareDiameter
0019|SIEMENS RA PLANE A|80|SS|1|CollimaterFingerTurnAngle
0019|SIEMENS RA PLANE A|82|SS|1|CollimaterFingerPosition
0019|SIEMENS RA PLANE A|84|SS|1|CollimaterDiaphragmTurnAngle
0019|SIEMENS RA PLANE A|86|SS|1|CollimaterDiaphragmPosition1
0019|SIEMENS RA PLANE A|88|SS|1|CollimaterDiaphragmPosition2
0019|SIEMENS RA PLANE A|8a|SS|1|CollimaterDiaphragmMode
0019|SIEMENS RA PLANE A|8c|SS|1|CollimaterBeamLimitBreadth
0019|SIEMENS RA PLANE A|8e|SS|1|CollimaterBeamLimitHeight
0019|SIEMENS RA PLANE A|90|SS|1|CollimaterBeamLimitDiameter
0019|SIEMENS RA PLANE A|92|SS|1|X-RayControlMOde
0019|SIEMENS RA PLANE A|94|SS|1|X-RaySystem
0019|SIEMENS RA PLANE A|96|SS|1|FocalSpot
0019|SIEMENS RA PLANE A|98|SS|1|ExposureControl
0019|SIEMENS RA PLANE A|9a|SL|1|XRayVoltage
0019|SIEMENS RA PLANE A|9c|SL|1|XRayCurrent
0019|SIEMENS RA PLANE A|9e|SL|1|XRayCurrentTimeProduct
0019|SIEMENS RA PLANE A|a0|SL|1|XRayPulseTime
0019|SIEMENS RA PLANE A|a2|SL|1|XRaySceneTimeFluoroClock
0019|SIEMENS RA PLANE A|a4|SS|1|MaximumPulseRate
0019|SIEMENS RA PLANE A|a6|SS|1|PulsesPerScene
0019|SIEMENS RA PLANE A|a8|SL|1|DoseAreaProductOfScene
0019|SIEMENS RA PLANE A|aa|SS|1|Dose
0019|SIEMENS RA PLANE A|ac|SS|1|DoseRate
0019|SIEMENS RA PLANE A|ae|SL|1|IIToCoverDistance
0019|SIEMENS RA PLANE A|b0|SS|1|LastFramePhase1
0019|SIEMENS RA PLANE A|b1|SS|1|FrameRatePhase1
0019|SIEMENS RA PLANE A|b2|SS|1|LastFramePhase2
0019|SIEMENS RA PLANE A|b3|SS|1|FrameRatePhase2
0019|SIEMENS RA PLANE A|b4|SS|1|LastFramePhase3
0019|SIEMENS RA PLANE A|b5|SS|1|FrameRatePhase3
0019|SIEMENS RA PLANE A|b6|SS|1|LastFramePhase4
0019|SIEMENS RA PLANE A|b7|SS|1|FrameRatePhase4
0019|SIEMENS RA PLANE A|b8|SS|1|GammaOfNativeImage
0019|SIEMENS RA PLANE A|b9|SS|1|GammaOfTVSystem
0019|SIEMENS RA PLANE A|bb|SL|1|PixelshiftX
0019|SIEMENS RA PLANE A|bc|SL|1|PixelshiftY
0019|SIEMENS RA PLANE A|bd|SL|1|MaskAverageFactor
0019|SIEMENS RA PLANE A|be|SL|1|BlankingCircleFlag
0019|SIEMENS RA PLANE A|bf|SL|1|CircleRowStart
0019|SIEMENS RA PLANE A|c0|SL|1|CircleRowEnd
0019|SIEMENS RA PLANE A|c1|SL|1|CircleColumnStart
0019|SIEMENS RA PLANE A|c2|SL|1|CircleColumnEnd
0019|SIEMENS RA PLANE A|c3|SL|1|CircleDiameter
0019|SIEMENS RA PLANE A|c4|SL|1|RectangularCollimaterFlag
0019|SIEMENS RA PLANE A|c5|SL|1|RectangleRowStart
0019|SVISION|90|LO|1|DeskCommand
0019|SIEMENS RA PLANE A|c6|SL|1|RectangleRowEnd
0019|SIEMENS RA PLANE A|c7|SL|1|RectangleColumnStart
0019|SIEMENS RA PLANE A|c8|SL|1|RectangleColumnEnd
0019|SIEMENS RA PLANE A|c9|SL|1|RectangleAngulation
0019|SIEMENS RA PLANE A|ca|SL|1|IrisCollimatorFlag
0019|SIEMENS RA PLANE A|cb|SL|1|IrisRowStart
0019|SIEMENS RA PLANE A|cc|SL|1|IrisRowEnd
0019|SIEMENS RA PLANE A|cd|SL|1|IrisColumnStart
0019|SIEMENS RA PLANE A|ce|SL|1|IrisColumnEnd
0019|SIEMENS RA PLANE A|cf|SL|1|IrisAngulation
0019|SIEMENS RA PLANE A|d1|SS|1|NumberOfFramesPlane
0019|SIEMENS RA PLANE A|d2|SS|1|Internal
0019|SIEMENS RA PLANE A|d3|SS|1|Internal
0019|SIEMENS RA PLANE A|d4|SS|1|Internal
0019|SIEMENS RA PLANE A|d5|SS|1|Internal
0019|SIEMENS RA PLANE A|d6|SS|1-n|Internal
0019|SIEMENS RA PLANE A|d7|SS|1-n|Internal
0019|SIEMENS RA PLANE A|d8|SS|1|Internal
0019|SIEMENS RA PLANE A|d9|SS|1|Internal
0019|SIEMENS RA PLANE A|da|SS|1|Internal
0019|SIEMENS RA PLANE A|db|SS|1|Internal
0019|SIEMENS RA PLANE A|dc|SS|1|Internal
0019|SIEMENS RA PLANE A|dd|SL|1|AnatomicBackground
0019|SIEMENS RA PLANE A|de|SL|1-n|AutoWindowBase
0019|SIEMENS RA PLANE A|df|SS|1|Internal
0019|SIEMENS RA PLANE A|e0|SL|1|Internal
0011|SIEMENS RA PLANE B|28|SL|1|FluoroTimerB
0011|SIEMENS RA PLANE B|29|SL|1|FluoroSkinDoseB
0011|SIEMENS RA PLANE B|2a|SL|1|TotalSkinDoseB
0011|SIEMENS RA PLANE B|2b|SL|1|FluoroDoseAreaProductB
0011|SIEMENS RA PLANE B|2c|SL|1|TotalDoseAreaProductB
0019|SIEMENS RA PLANE B|18|SS|1|Internal
0019|SIEMENS RA PLANE B|19|SS|1|Internal
0019|SIEMENS RA PLANE B|1a|SS|1|Internal
0019|SIEMENS RA PLANE B|1b|SS|1|Internal
0019|SIEMENS RA PLANE B|1c|SS|1|Internal
0019|SIEMENS RA PLANE B|1d|SS|1|Internal
0019|SIEMENS RA PLANE B|1e|SS|1|Internal
0019|SIEMENS RA PLANE B|1f|SS|1|Internal
0019|SIEMENS RA PLANE B|20|SL|1-n|SystemCalibFactorPlaneB
0019|SIEMENS RA PLANE B|22|US|1|Unknown
0019|SIEMENS RA PLANE B|24|US|1|Unknown
0019|SIEMENS RA PLANE B|26|US|1|Unknown
0019|SIEMENS RA PLANE B|28|US|1|Unknown
0019|SIEMENS RA PLANE B|2a|US|1|Unknown
0019|SIEMENS RA PLANE B|2c|US|1|Unknown
0019|SIEMENS RA PLANE B|2e|US|1|Unknown
0019|SIEMENS RA PLANE B|30|US|1|Unknown
0019|SIEMENS RA PLANE B|32|US|1|Unknown
0019|SIEMENS RA PLANE B|34|US|1|Unknown
0019|SIEMENS RA PLANE B|36|US|1|Unknown
0019|SIEMENS RA PLANE B|38|US|1|Unknown
0019|SIEMENS RA PLANE B|3a|US|1|Unknown
0019|SIEMENS RA PLANE B|3c|US|1|Unknown
0019|SIEMENS RA PLANE B|3e|US|1|Unknown
0019|SIEMENS RA PLANE B|40|US|1|Unknown
0019|SIEMENS RA PLANE B|42|US|1|Unknown
0019|SIEMENS RA PLANE B|44|US|1|Unknown
0019|SIEMENS RA PLANE B|46|US|1|Unknown
0019|SIEMENS RA PLANE B|48|US|1|Unknown
0019|SIEMENS RA PLANE B|4a|US|1-n|Unknown
0019|SIEMENS RA PLANE B|4c|US|1-n|Unknown
0019|SIEMENS RA PLANE B|4e|US|1-n|Unknown
0019|SIEMENS RA PLANE B|50|US|1|Unknown
0019|SIEMENS RA PLANE B|52|US|1|Unknown
0019|SIEMENS RA PLANE B|54|US|1|Unknown
0019|SIEMENS RA PLANE B|56|US|1|Unknown
0019|SIEMENS RA PLANE B|58|US|1|Unknown
0019|SIEMENS RA PLANE B|5a|US|1|Unknown
0019|SIEMENS RA PLANE B|5c|US|1-n|Unknown
0019|SIEMENS RA PLANE B|5e|US|1-n|Unknown
0019|SIEMENS RA PLANE B|60|US|1-n|Unknown
0019|SIEMENS RA PLANE B|62|US|1-n|Unknown
0019|SIEMENS RA PLANE B|64|US|1-n|Unknown
0019|SIEMENS RA PLANE B|66|US|1-n|Unknown
0019|SIEMENS RA PLANE B|68|US|1-n|Unknown
0019|SIEMENS RA PLANE B|6a|US|1-n|Unknown
0019|SIEMENS RA PLANE B|6c|US|1-n|Unknown
0019|SIEMENS RA PLANE B|6e|US|1-n|Unknown
0019|SIEMENS RA PLANE B|70|US|1-n|Unknown
0019|SIEMENS RA PLANE B|72|UN|1|Unknown
0019|SIEMENS RA PLANE B|74|UN|1|Unknown
0019|SIEMENS RA PLANE B|76|UN|1|Unknown
0019|SIEMENS RA PLANE B|78|US|1-n|Unknown
0019|SIEMENS RA PLANE B|7a|US|1|Unknown
0019|SIEMENS RA PLANE B|7c|US|1|Unknown
0019|SIEMENS RA PLANE B|7e|US|1|Unknown
0019|SIEMENS RA PLANE B|80|US|1|Unknown
0019|SIEMENS RA PLANE B|82|US|1|Unknown
0019|SIEMENS RA PLANE B|84|US|1|Unknown
0019|SIEMENS RA PLANE B|86|US|1|Unknown
0019|SIEMENS RA PLANE B|88|US|1|Unknown
0019|SIEMENS RA PLANE B|8a|US|1|Unknown
0019|SIEMENS RA PLANE B|8c|US|1|Unknown
0019|SIEMENS RA PLANE B|8e|US|1|Unknown
0019|SIEMENS RA PLANE B|90|US|1|Unknown
0019|SIEMENS RA PLANE B|92|US|1|Unknown
0019|SIEMENS RA PLANE B|94|US|1|Unknown
0019|SIEMENS RA PLANE B|96|US|1|Unknown
0019|SIEMENS RA PLANE B|98|US|1|Unknown
0019|SIEMENS RA PLANE B|9a|US|1-n|Unknown
0019|SIEMENS RA PLANE B|9c|US|1-n|Unknown
0019|SIEMENS RA PLANE B|9e|US|1-n|Unknown
0019|SIEMENS RA PLANE B|a0|US|1-n|Unknown
0019|SIEMENS RA PLANE B|a2|US|1-n|Unknown
0019|SIEMENS RA PLANE B|a4|US|1|Unknown
0019|SIEMENS RA PLANE B|a6|US|1|Unknown
0019|SIEMENS RA PLANE B|a8|US|1-n|Unknown
0019|SIEMENS RA PLANE B|aa|US|1|Unknown
0019|SIEMENS RA PLANE B|ac|US|1|Unknown
0011|SIEMENS RIS|10|LT|1|PatientUID
0011|SIEMENS RIS|11|LT|1|PatientID
0011|SIEMENS RIS|20|DA|1|PatientRegistrationDate
0011|SIEMENS RIS|21|TM|1|PatientRegistrationTime
0011|SIEMENS RIS|30|LT|1|PatientnameRIS
0011|SIEMENS RIS|31|LT|1|PatientprenameRIS
0011|SIEMENS RIS|40|LT|1|PatientHospitalStatus
0011|SIEMENS RIS|41|LT|1|MedicalAlerts
0011|SIEMENS RIS|42|LT|1|ContrastAllergies
0031|SIEMENS RIS|10|LT|1|RequestUID
0031|SIEMENS RIS|45|LT|1|RequestingPhysician
0031|SIEMENS RIS|50|LT|1|RequestedPhysician
0033|SIEMENS RIS|10|LT|1|PatientStudyUID
0021|SIEMENS SMS-AX  ACQ 1.0|00|US|1|AcquisitionType
0021|SIEMENS SMS-AX  ACQ 1.0|01|US|1|AcquisitionMode
0021|SIEMENS SMS-AX  ACQ 1.0|02|US|1|FootswitchIndex
0021|SIEMENS SMS-AX  ACQ 1.0|03|US|1|AcquisitionRoom
0021|SIEMENS SMS-AX  ACQ 1.0|04|SL|1|CurrentTimeProduct
0021|SIEMENS SMS-AX  ACQ 1.0|05|SL|1|Dose
0021|SIEMENS SMS-AX  ACQ 1.0|06|SL|1|SkinDosePercent
0021|SIEMENS SMS-AX  ACQ 1.0|07|SL|1|SkinDoseAccumulation
0021|SIEMENS SMS-AX  ACQ 1.0|08|SL|1|SkinDoseRate
0021|SIEMENS SMS-AX  ACQ 1.0|0A|UL|1|CopperFilter
0021|SIEMENS SMS-AX  ACQ 1.0|0B|US|1|MeasuringField
0021|SIEMENS SMS-AX  ACQ 1.0|0C|SS|3|PostBlankingCircle
0021|SIEMENS SMS-AX  ACQ 1.0|0D|SS|2-2n|DynaAngles
0021|SIEMENS SMS-AX  ACQ 1.0|0E|SS|1|TotalSteps
0021|SIEMENS SMS-AX  ACQ 1.0|0F|SL|3-3n|DynaXRayInfo
0021|SIEMENS SMS-AX  ACQ 1.0|10|US|1|ModalityLUTInputGamma
0021|SIEMENS SMS-AX  ACQ 1.0|11|US|1|ModalityLUTOutputGamma
0021|SIEMENS SMS-AX  ACQ 1.0|12|OB|1-n|SH_STPAR
0021|SIEMENS SMS-AX  ACQ 1.0|13|US|1|AcquisitionZoom
0021|SIEMENS SMS-AX  ACQ 1.0|14|SS|1|DynaAngulationStepWidth
0021|SIEMENS SMS-AX  ACQ 1.0|15|US|1|Harmonization
0021|SIEMENS SMS-AX  ACQ 1.0|16|US|1|DRSingleFlag
0021|SIEMENS SMS-AX  ACQ 1.0|17|SL|1|SourceToIsocenter
0021|SIEMENS SMS-AX  ACQ 1.0|18|US|1|PressureData
0021|SIEMENS SMS-AX  ACQ 1.0|19|SL|1|ECGIndexArray
0021|SIEMENS SMS-AX  ACQ 1.0|1A|US|1|FDFlag
0021|SIEMENS SMS-AX  ACQ 1.0|1B|OB|1|SH_ZOOM
0021|SIEMENS SMS-AX  ACQ 1.0|1C|OB|1|SH_COLPAR
0021|SIEMENS SMS-AX  ACQ 1.0|1D|US|1|K_Factor
0021|SIEMENS SMS-AX  ACQ 1.0|1E|US|8|EVE
0021|SIEMENS SMS-AX  ACQ 1.0|1F|SL|1|TotalSceneTime
0021|SIEMENS SMS-AX  ACQ 1.0|20|US|1|RestoreFlag
0021|SIEMENS SMS-AX  ACQ 1.0|21|US|1|StandMovementFlag
0021|SIEMENS SMS-AX  ACQ 1.0|22|US|1|FDRows
0021|SIEMENS SMS-AX  ACQ 1.0|23|US|1|FDColumns
0021|SIEMENS SMS-AX  ACQ 1.0|24|US|1|TableMovementFlag
0021|SIEMENS SMS-AX  ACQ 1.0|25|LO|1|OriginalOrganProgramName
0021|SIEMENS SMS-AX  ACQ 1.0|26|DS|1|CrispyXPIFilter
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|00|US|1|ViewNative
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|01|US|1|OriginalSeriesNumber
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|02|US|1|OriginalImageNumber
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|03|US|1|WinCenter
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|04|US|1|WinWidth
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|05|US|1|WinBrightness
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|06|US|1|WinContrast
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|07|US|1|OriginalFrameNumber
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|08|US|1|OriginalMaskFrameNumber
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|09|US|1|Opac
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0A|US|1|OriginalNumberOfFrames
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0B|DS|1|OriginalSceneDuration
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0C|LO|1|IdentifierLOID
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0D|SS|1-n|OriginalSceneVFRInfo
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0E|SS|1|OriginalFrameECGPosition
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0F|SS|1|OriginalECG1stFrameOffset_retired
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|10|SS|1|ZoomFlag
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|11|US|1|Flex
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|12|US|1|NumberOfMaskFrames
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|13|US|1|NumberOfFillFrames
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|14|US|1|SeriesNumber
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|15|IS|1|ImageNumber
0023|SIEMENS SMS-AX  QUANT 1.0|00|DS|2|HorizontalCalibrationPixelSize
0023|SIEMENS SMS-AX  QUANT 1.0|01|DS|2|VerticalCalibrationPixelSize
0023|SIEMENS SMS-AX  QUANT 1.0|02|LO|1|CalibrationObject
0023|SIEMENS SMS-AX  QUANT 1.0|03|DS|1|CalibrationObjectSize
0023|SIEMENS SMS-AX  QUANT 1.0|04|LO|1|CalibrationMethod
0023|SIEMENS SMS-AX  QUANT 1.0|05|ST|1|Filename
0023|SIEMENS SMS-AX  QUANT 1.0|06|IS|1|FrameNumber
0023|SIEMENS SMS-AX  QUANT 1.0|07|IS|2|CalibrationFactorMultiplicity
0023|SIEMENS SMS-AX  QUANT 1.0|08|IS|1|CalibrationTODValue
0019|SIEMENS SMS-AX  VIEW 1.0|00|US|1|ReviewMode
0019|SIEMENS SMS-AX  VIEW 1.0|01|US|1|AnatomicalBackgroundPercent
0019|SIEMENS SMS-AX  VIEW 1.0|02|US|1|NumberOfPhases
0019|SIEMENS SMS-AX  VIEW 1.0|03|US|1|ApplyAnatomicalBackground
0019|SIEMENS SMS-AX  VIEW 1.0|04|SS|4-4n|PixelShiftArray
0019|SIEMENS SMS-AX  VIEW 1.0|05|US|1|Brightness
0019|SIEMENS SMS-AX  VIEW 1.0|06|US|1|Contrast
0019|SIEMENS SMS-AX  VIEW 1.0|07|US|1|Enabled
0019|SIEMENS SMS-AX  VIEW 1.0|08|US|1|NativeEdgeEnhancementPercentGain
0019|SIEMENS SMS-AX  VIEW 1.0|09|SS|1|NativeEdgeEnhancementLUTIndex
0019|SIEMENS SMS-AX  VIEW 1.0|0A|SS|1|NativeEdgeEnhancementKernelSize
0019|SIEMENS SMS-AX  VIEW 1.0|0B|US|1|SubtrEdgeEnhancementPercentGain
0019|SIEMENS SMS-AX  VIEW 1.0|0C|SS|1|SubtrEdgeEnhancementLUTIndex
0019|SIEMENS SMS-AX  VIEW 1.0|0D|SS|1|SubtrEdgeEnhancementKernelSize
0019|SIEMENS SMS-AX  VIEW 1.0|0E|US|1|FadePercent
0019|SIEMENS SMS-AX  VIEW 1.0|0F|US|1|FlippedBeforeLateralityApplied
0019|SIEMENS SMS-AX  VIEW 1.0|10|US|1|ApplyFade
0019|SIEMENS SMS-AX  VIEW 1.0|12|US|1|Zoom
0019|SIEMENS SMS-AX  VIEW 1.0|13|SS|1|PanX
0019|SIEMENS SMS-AX  VIEW 1.0|14|SS|1|PanY
0019|SIEMENS SMS-AX  VIEW 1.0|15|SS|1|NativeEdgeEnhancementAdvPercGain
0019|SIEMENS SMS-AX  VIEW 1.0|16|SS|1|SubtrEdgeEnhancementAdvPercGain
0019|SIEMENS SMS-AX  VIEW 1.0|17|US|1|InvertFlag
0019|SIEMENS SMS-AX  VIEW 1.0|1A|OB|1|Quant1KOverlay
0019|SIEMENS SMS-AX  VIEW 1.0|1B|US|1|OriginalResolution
0019|SIEMENS SMS-AX  VIEW 1.0|1C|DS|1|AutoWindowCenter
0019|SIEMENS SMS-AX  VIEW 1.0|1D|DS|1|AutoWindowWidth
0009|SIENET|01|US|1|SIENETCommandField
0009|SIENET|14|LT|1|ReceiverPLA
0009|SIENET|16|US|1|TransferPriority
0009|SIENET|29|LT|1|ActualUser
0095|SIENET|01|LT|1|ExaminationFolderID
0095|SIENET|04|UL|1|FolderReportedStatus
0095|SIENET|05|LT|1|FolderReportingRadiologist
0095|SIENET|07|LT|1|SIENETISAPLA
0099|SIENET|02|UL|1|DataObjectAttributes
0009|SPI RELEASE 1|10|LT|1|Comments
0009|SPI RELEASE 1|15|LO|1|SPIImageUID
0009|SPI RELEASE 1|40|US|1|DataObjectType
0009|SPI RELEASE 1|41|LO|1|DataObjectSubtype
0011|SPI RELEASE 1|10|LO|1|Organ
0011|SPI RELEASE 1|15|LO|1|AllergyIndication
0011|SPI RELEASE 1|20|LO|1|Pregnancy
0029|SPI RELEASE 1|60|LT|1|CompressionAlgorithm
0009|SPI Release 1|10|LT|1|Comments
0009|SPI Release 1|15|LO|1|SPIImageUID
0009|SPI Release 1|40|US|1|DataObjectType
0009|SPI Release 1|41|LO|1|DataObjectSubtype
0011|SPI Release 1|10|LO|1|Organ
0011|SPI Release 1|15|LO|1|AllergyIndication
0011|SPI Release 1|20|LO|1|Pregnancy
0029|SPI Release 1|60|LT|1|CompressionAlgorithm
0009|SPI|10|LO|1|Comments
0009|SPI|15|LO|1|SPIImageUID
0009|SPI|40|US|1|DataObjectType
0009|SPI|41|LT|1|DataObjectSubtype
0011|SPI|10|LT|1|Organ
0011|SPI|15|LT|1|AllergyIndication
0011|SPI|20|LT|1|Pregnancy
0029|SPI|60|LT|1|CompressionAlgorithm
0009|SPI-P Release 1|00|LT|1|DataObjectRecognitionCode
0009|SPI-P Release 1|04|LO|1|ImageDataConsistence
0009|SPI-P Release 1|08|US|1|Unknown
0009|SPI-P Release 1|12|LO|1|Unknown
0009|SPI-P Release 1|15|LO|1|UniqueIdentifier
0009|SPI-P Release 1|16|LO|1|Unknown
0009|SPI-P Release 1|18|LO|1|Unknown
0009|SPI-P Release 1|21|LT|1|Unknown
0009|SPI-P Release 1|31|LT|1|PACSUniqueIdentifier
0009|SPI-P Release 1|34|LT|1|ClusterUniqueIdentifier
0009|SPI-P Release 1|38|LT|1|SystemUniqueIdentifier
0009|SPI-P Release 1|39|LT|1|Unknown
0009|SPI-P Release 1|51|LT|1|StudyUniqueIdentifier
0009|SPI-P Release 1|61|LT|1|SeriesUniqueIdentifier
0009|SPI-P Release 1|91|LT|1|Unknown
0009|SPI-P Release 1|f2|LT|1|Unknown
0009|SPI-P Release 1|f3|UN|1|Unknown
0009|SPI-P Release 1|f4|LT|1|Unknown
0009|SPI-P Release 1|f5|UN|1|Unknown
0009|SPI-P Release 1|f7|LT|1|Unknown
0011|SPI-P Release 1|10|LT|1|PatientEntryID
0011|SPI-P Release 1|21|UN|1|Unknown
0011|SPI-P Release 1|22|UN|1|Unknown
0011|SPI-P Release 1|31|UN|1|Unknown
0011|SPI-P Release 1|32|UN|1|Unknown
0019|SPI-P Release 1|00|UN|1|Unknown
0019|SPI-P Release 1|01|UN|1|Unknown
0019|SPI-P Release 1|02|UN|1|Unknown
0019|SPI-P Release 1|10|US|1|MainsFrequency
0019|SPI-P Release 1|25|LT|1-n|OriginalPixelDataQuality
0019|SPI-P Release 1|30|US|1|ECGTriggering
0019|SPI-P Release 1|31|UN|1|ECG1Offset
0019|SPI-P Release 1|32|UN|1|ECG2Offset1
0019|SPI-P Release 1|33|UN|1|ECG2Offset2
0019|SPI-P Release 1|50|US|1|VideoScanMode
0019|SPI-P Release 1|51|US|1|VideoLineRate
0019|SPI-P Release 1|60|US|1|XrayTechnique
0019|SPI-P Release 1|61|DS|1|ImageIdentifierFromat
0019|SPI-P Release 1|62|US|1|IrisDiaphragm
0019|SPI-P Release 1|63|CS|1|Filter
0019|SPI-P Release 1|64|CS|1|CineParallel
0019|SPI-P Release 1|65|CS|1|CineMaster
0019|SPI-P Release 1|70|US|1|ExposureChannel
0019|SPI-P Release 1|71|UN|1|ExposureChannelFirstImage
0019|SPI-P Release 1|72|US|1|ProcessingChannel
0019|SPI-P Release 1|80|DS|1|AcquisitionDelay
0019|SPI-P Release 1|81|UN|1|RelativeImageTime
0019|SPI-P Release 1|90|CS|1|VideoWhiteCompression
0019|SPI-P Release 1|a0|US|1|Angulation
0019|SPI-P Release 1|a1|US|1|Rotation
0021|SPI-P Release 1|12|LT|1|SeriesUniqueIdentifier
0021|SPI-P Release 1|14|LT|1|Unknown
0029|SPI-P Release 1|00|DS|4|Unknown
0029|SPI-P Release 1|20|DS|1|PixelAspectRatio
0029|SPI-P Release 1|25|LO|1-n|ProcessedPixelDataQuality
0029|SPI-P Release 1|30|LT|1|Unknown
0029|SPI-P Release 1|38|US|1|Unknown
0029|SPI-P Release 1|60|LT|1|Unknown
0029|SPI-P Release 1|61|LT|1|Unknown
0029|SPI-P Release 1|67|LT|1|Unknown
0029|SPI-P Release 1|70|LT|1|WindowID
0029|SPI-P Release 1|71|CS|1|VideoInvertSubtracted
0029|SPI-P Release 1|72|CS|1|VideoInvertNonsubtracted
0029|SPI-P Release 1|77|CS|1|WindowSelectStatus
0029|SPI-P Release 1|78|LT|1|ECGDisplayPrintingID
0029|SPI-P Release 1|79|CS|1|ECGDisplayPrinting
0029|SPI-P Release 1|7e|CS|1|ECGDisplayPrintingEnableStatus
0029|SPI-P Release 1|7f|CS|1|ECGDisplayPrintingSelectStatus
0029|SPI-P Release 1|80|LT|1|PhysiologicalDisplayID
0029|SPI-P Release 1|81|US|1|PreferredPhysiologicalChannelDisplay
0029|SPI-P Release 1|8e|CS|1|PhysiologicalDisplayEnableStatus
0029|SPI-P Release 1|8f|CS|1|PhysiologicalDisplaySelectStatus
0029|SPI-P Release 1|c0|LT|1|FunctionalShutterID
0029|SPI-P Release 1|c1|US|1|FieldOfShutter
0029|SPI-P Release 1|c5|LT|1|FieldOfShutterRectangle
0029|SPI-P Release 1|ce|CS|1|ShutterEnableStatus
0029|SPI-P Release 1|cf|CS|1|ShutterSelectStatus
7FE1|SPI-P Release 1|10|ox|1|PixelData
0009|SPI-P Release 1;1|c0|LT|1|Unknown
0009|SPI-P Release 1;1|c1|LT|1|Unknown
0019|SPI-P Release 1;1|00|UN|1|PhysiologicalDataType
0019|SPI-P Release 1;1|01|UN|1|PhysiologicalDataChannelAndKind
0019|SPI-P Release 1;1|02|US|1|SampleBitsAllocated
0019|SPI-P Release 1;1|03|US|1|SampleBitsStored
0019|SPI-P Release 1;1|04|US|1|SampleHighBit
0019|SPI-P Release 1;1|05|US|1|SampleRepresentation
0019|SPI-P Release 1;1|06|UN|1|SmallestSampleValue
0019|SPI-P Release 1;1|07|UN|1|LargestSampleValue
0019|SPI-P Release 1;1|08|UN|1|NumberOfSamples
0019|SPI-P Release 1;1|09|UN|1|SampleData
0019|SPI-P Release 1;1|0a|UN|1|SampleRate
0019|SPI-P Release 1;1|10|UN|1|PhysiologicalDataType2
0019|SPI-P Release 1;1|11|UN|1|PhysiologicalDataChannelAndKind2
0019|SPI-P Release 1;1|12|US|1|SampleBitsAllocated2
0019|SPI-P Release 1;1|13|US|1|SampleBitsStored2
0019|SPI-P Release 1;1|14|US|1|SampleHighBit2
0019|SPI-P Release 1;1|15|US|1|SampleRepresentation2
0019|SPI-P Release 1;1|16|UN|1|SmallestSampleValue2
0019|SPI-P Release 1;1|17|UN|1|LargestSampleValue2
0019|SPI-P Release 1;1|18|UN|1|NumberOfSamples2
0019|SPI-P Release 1;1|19|UN|1|SampleData2
0019|SPI-P Release 1;1|1a|UN|1|SampleRate2
0029|SPI-P Release 1;1|00|LT|1|ZoomID
0029|SPI-P Release 1;1|01|DS|1-n|ZoomRectangle
0029|SPI-P Release 1;1|03|DS|1|ZoomFactor
0029|SPI-P Release 1;1|04|US|1|ZoomFunction
0029|SPI-P Release 1;1|0e|CS|1|ZoomEnableStatus
0029|SPI-P Release 1;1|0f|CS|1|ZoomSelectStatus
0029|SPI-P Release 1;1|40|LT|1|MagnifyingGlassID
0029|SPI-P Release 1;1|41|DS|1-n|MagnifyingGlassRectangle
0029|SPI-P Release 1;1|43|DS|1|MagnifyingGlassFactor
0029|SPI-P Release 1;1|44|US|1|MagnifyingGlassFunction
0029|SPI-P Release 1;1|4e|CS|1|MagnifyingGlassEnableStatus
0029|SPI-P Release 1;1|4f|CS|1|MagnifyingGlassSelectStatus
0029|SPI-P Release 1;2|00|LT|1|SubtractionMaskID
0029|SPI-P Release 1;2|04|UN|1|MaskingFunction
0029|SPI-P Release 1;2|0c|UN|1|ProprietaryMaskingParameters
0029|SPI-P Release 1;2|1e|CS|1|SubtractionMaskEnableStatus
0029|SPI-P Release 1;2|1f|CS|1|SubtractionMaskSelectStatus
0029|SPI-P Release 1;3|00|LT|1|ImageEnhancementID
0029|SPI-P Release 1;3|01|LT|1|ImageEnhancement
0029|SPI-P Release 1;3|02|LT|1|ConvolutionID
0029|SPI-P Release 1;3|03|LT|1|ConvolutionType
0029|SPI-P Release 1;3|04|LT|1|ConvolutionKernelSizeID
0029|SPI-P Release 1;3|05|US|2|ConvolutionKernelSize
0029|SPI-P Release 1;3|06|US|1-n|ConvolutionKernel
0029|SPI-P Release 1;3|0c|DS|1|EnhancementGain
0029|SPI-P Release 1;3|1e|CS|1|ImageEnhancementEnableStatus
0029|SPI-P Release 1;3|1f|CS|1|ImageEnhancementSelectStatus
0011|SPI-P Release 2;1|18|LT|1|Unknown
0023|SPI-P Release 2;1|0d|UI|1|Unknown
0023|SPI-P Release 2;1|0e|UI|1|Unknown
0009|SPI-P-GV-CT Release 1|00|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|10|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|20|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|30|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|40|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|50|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|60|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|70|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|75|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|80|LO|1|Unknown
0009|SPI-P-GV-CT Release 1|90|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|08|IS|1|Unknown
0019|SPI-P-GV-CT Release 1|09|IS|1|Unknown
0019|SPI-P-GV-CT Release 1|0a|IS|1|Unknown
0019|SPI-P-GV-CT Release 1|10|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|20|TM|1|Unknown
0019|SPI-P-GV-CT Release 1|50|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|60|DS|1|Unknown
0019|SPI-P-GV-CT Release 1|61|US|1|Unknown
0019|SPI-P-GV-CT Release 1|63|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|64|US|1|Unknown
0019|SPI-P-GV-CT Release 1|65|IS|1|Unknown
0019|SPI-P-GV-CT Release 1|70|LT|1|Unknown
0019|SPI-P-GV-CT Release 1|80|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|81|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|90|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|a0|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|a1|US|1|Unknown
0019|SPI-P-GV-CT Release 1|a2|US|1|Unknown
0019|SPI-P-GV-CT Release 1|a3|US|1|Unknown
0019|SPI-P-GV-CT Release 1|b0|LO|1|Unknown
0019|SPI-P-GV-CT Release 1|b1|LO|1|Unknown
0021|SPI-P-GV-CT Release 1|20|LO|1|Unknown
0021|SPI-P-GV-CT Release 1|30|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|40|LO|1|Unknown
0021|SPI-P-GV-CT Release 1|50|LO|1|Unknown
0021|SPI-P-GV-CT Release 1|60|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|70|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|80|DS|1|Unknown
0019|SVISION|A0|DS|1|ExtendedExposureTime
0021|SPI-P-GV-CT Release 1|90|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|a0|US|1|Unknown
0021|SPI-P-GV-CT Release 1|a1|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|a2|DS|1|Unknown
0021|SPI-P-GV-CT Release 1|a3|LT|1|Unknown
0021|SPI-P-GV-CT Release 1|a4|LT|1|Unknown
0021|SPI-P-GV-CT Release 1|b0|LO|1|Unknown
0021|SPI-P-GV-CT Release 1|c0|LO|1|Unknown
0029|SPI-P-GV-CT Release 1|10|LO|1|Unknown
0029|SPI-P-GV-CT Release 1|30|UL|1|Unknown
0029|SPI-P-GV-CT Release 1|31|UL|1|Unknown
0029|SPI-P-GV-CT Release 1|32|UL|1|Unknown
0029|SPI-P-GV-CT Release 1|33|UL|1|Unknown
0029|SPI-P-GV-CT Release 1|80|LO|1|Unknown
0029|SPI-P-GV-CT Release 1|90|LO|1|Unknown
0029|SPI-P-GV-CT Release 1|d0|IS|1|Unknown
0029|SPI-P-GV-CT Release 1|d1|IS|1|Unknown
0019|SPI-P-PCR Release 2|30|US|1|Unknown
0021|SPI-P-Private-CWS Release 1|00|LT|1|WindowOfImagesID
0021|SPI-P-Private-CWS Release 1|01|CS|1|WindowOfImagesType
0021|SPI-P-Private-CWS Release 1|02|IS|1-n|WindowOfImagesScope
0019|SPI-P-Private-DCI Release 1|10|UN|1|ECGTimeMapDataBitsAllocated
0019|SPI-P-Private-DCI Release 1|11|UN|1|ECGTimeMapDataBitsStored
0019|SPI-P-Private-DCI Release 1|12|UN|1|ECGTimeMapDataHighBit
0019|SPI-P-Private-DCI Release 1|13|UN|1|ECGTimeMapDataRepresentation
0019|SPI-P-Private-DCI Release 1|14|UN|1|ECGTimeMapDataSmallestDataValue
0019|SPI-P-Private-DCI Release 1|15|UN|1|ECGTimeMapDataLargestDataValue
0019|SPI-P-Private-DCI Release 1|16|UN|1|ECGTimeMapDataNumberOfDataValues
0019|SPI-P-Private-DCI Release 1|17|UN|1|ECGTimeMapData
0021|SPI-P-Private_CDS Release 1|40|IS|1|Unknown
0029|SPI-P-Private_CDS Release 1|00|UN|1|Unknown
0019|SPI-P-Private_ICS Release 1|30|DS|1|Unknown
0019|SPI-P-Private_ICS Release 1|31|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1|08|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|0f|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|10|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|1b|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|1c|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|21|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|43|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|44|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|4C|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|67|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1|68|US|1|Unknown
0029|SPI-P-Private_ICS Release 1|6A|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1|6B|US|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|00|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|05|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|06|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|20|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|21|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|CD|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|00|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|01|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|02|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|03|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|04|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|05|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C0|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C1|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C2|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C3|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C4|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|C5|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|02|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|9A|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|E0|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;5|50|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1;5|55|CS|1|Unknown
0019|SPI-P-XSB-DCI Release 1|10|LT|1|VideoBeamBoost
0019|SPI-P-XSB-DCI Release 1|11|US|1|ChannelGeneratingVideoSync
0019|SPI-P-XSB-DCI Release 1|12|US|1|VideoGain
0019|SPI-P-XSB-DCI Release 1|13|US|1|VideoOffset
0019|SPI-P-XSB-DCI Release 1|20|DS|1|RTDDataCompressionFactor
0029|Silhouette Annot V1.0|11|IS|1|AnnotationName
0029|Silhouette Annot V1.0|12|LT|1|AnnotationFont
0029|Silhouette Annot V1.0|13|LT|1|AnnotationTextForegroundColor
0029|Silhouette Annot V1.0|14|LT|1|AnnotationTextBackgroundColor
0029|Silhouette Annot V1.0|15|UL|1|AnnotationTextBackingMode
0029|Silhouette Annot V1.0|16|UL|1|AnnotationTextJustification
0029|Silhouette Annot V1.0|17|UL|1|AnnotationTextLocation
0029|Silhouette Annot V1.0|18|LT|1|AnnotationTextString
0029|Silhouette Annot V1.0|19|UL|1|AnnotationTextAttachMode
0029|Silhouette Annot V1.0|20|UL|1|AnnotationTextCursorMode
0029|Silhouette Annot V1.0|21|UL|1|AnnotationTextShadowOffsetX
0029|Silhouette Annot V1.0|22|UL|1|AnnotationTextShadowOffsetY
0029|Silhouette Annot V1.0|23|LT|1|AnnotationLineColor
0029|Silhouette Annot V1.0|24|UL|1|AnnotationLineThickness
0029|Silhouette Annot V1.0|25|UL|1|AnnotationLineType
0029|Silhouette Annot V1.0|26|UL|1|AnnotationLineStyle
0029|Silhouette Annot V1.0|27|UL|1|AnnotationLineDashLength
0029|Silhouette Annot V1.0|28|UL|1|AnnotationLineAttachMode
0029|Silhouette Annot V1.0|29|UL|1|AnnotationLinePointCount
0029|Silhouette Annot V1.0|30|FD|1|AnnotationLinePoints
0019|SVISION|A1|DS|1|ActualExposureTime
0029|Silhouette Annot V1.0|31|UL|1|AnnotationLineControlSize
0029|Silhouette Annot V1.0|32|LT|1|AnnotationMarkerColor
0029|Silhouette Annot V1.0|33|UL|1|AnnotationMarkerType
0029|Silhouette Annot V1.0|34|UL|1|AnnotationMarkerSize
0029|Silhouette Annot V1.0|35|FD|1|AnnotationMarkerLocation
0029|Silhouette Annot V1.0|36|UL|1|AnnotationMarkerAttachMode
0029|Silhouette Annot V1.0|37|LT|1|AnnotationGeomColor
0029|Silhouette Annot V1.0|38|UL|1|AnnotationGeomThickness
0029|Silhouette Annot V1.0|39|UL|1|AnnotationGeomLineStyle
0029|Silhouette Annot V1.0|40|UL|1|AnnotationGeomDashLength
0029|Silhouette Annot V1.0|41|UL|1|AnnotationGeomFillPattern
0029|Silhouette Annot V1.0|42|UL|1|AnnotationInteractivity
0029|Silhouette Annot V1.0|43|FD|1|AnnotationArrowLength
0029|Silhouette Annot V1.0|44|FD|1|AnnotationArrowAngle
0029|Silhouette Annot V1.0|45|UL|1|AnnotationDontSave
0029|Silhouette Graphics Export V1.0|00|UI|1|Unknown
0029|Silhouette Line V1.0|11|IS|1|LineName
0029|Silhouette Line V1.0|12|LT|1|LineNameFont
0029|Silhouette Line V1.0|13|UL|1|LineNameDisplay
0029|Silhouette Line V1.0|14|LT|1|LineNormalColor
0029|Silhouette Line V1.0|15|UL|1|LineType
0029|Silhouette Line V1.0|16|UL|1|LineThickness
0029|Silhouette Line V1.0|17|UL|1|LineStyle
0029|Silhouette Line V1.0|18|UL|1|LineDashLength
0029|Silhouette Line V1.0|19|UL|1|LineInteractivity
0029|Silhouette Line V1.0|20|LT|1|LineMeasurementColor
0029|Silhouette Line V1.0|21|LT|1|LineMeasurementFont
0029|Silhouette Line V1.0|22|UL|1|LineMeasurementDashLength
0029|Silhouette Line V1.0|23|UL|1|LinePointSpace
0029|Silhouette Line V1.0|24|FD|1|LinePoints
0029|Silhouette Line V1.0|25|UL|1|LineControlPointSize
0029|Silhouette Line V1.0|26|UL|1|LineControlPointSpace
0029|Silhouette Line V1.0|27|FD|1|LineControlPoints
0029|Silhouette Line V1.0|28|LT|1|LineLabel
0029|Silhouette Line V1.0|29|UL|1|LineDontSave
0029|Silhouette ROI V1.0|11|IS|1|ROIName
0029|Silhouette ROI V1.0|12|LT|1|ROINameFont
0029|Silhouette ROI V1.0|13|LT|1|ROINormalColor
0029|Silhouette ROI V1.0|14|UL|1|ROIFillPattern
0029|Silhouette ROI V1.0|15|UL|1|ROIBpSeg
0029|Silhouette ROI V1.0|16|UN|1|ROIBpSegPairs
0029|Silhouette ROI V1.0|17|UL|1|ROISeedSpace
0029|Silhouette ROI V1.0|18|UN|1|ROISeeds
0029|Silhouette ROI V1.0|19|UL|1|ROILineThickness
0029|Silhouette ROI V1.0|20|UL|1|ROILineStyle
0029|Silhouette ROI V1.0|21|UL|1|ROILineDashLength
0029|Silhouette ROI V1.0|22|UL|1|ROIInteractivity
0029|Silhouette ROI V1.0|23|UL|1|ROINamePosition
0029|Silhouette ROI V1.0|24|UL|1|ROINameDisplay
0029|Silhouette ROI V1.0|25|LT|1|ROILabel
0029|Silhouette ROI V1.0|26|UL|1|ROIShape
0029|Silhouette ROI V1.0|27|FD|1|ROIShapeTilt
0029|Silhouette ROI V1.0|28|UL|1|ROIShapePointsCount
0029|Silhouette ROI V1.0|29|UL|1|ROIShapePointsSpace
0029|Silhouette ROI V1.0|30|FD|1|ROIShapePoints
0029|Silhouette ROI V1.0|31|UL|1|ROIShapeControlPointsCount
0029|Silhouette ROI V1.0|32|UL|1|ROIShapeControlPointsSpace
0029|Silhouette ROI V1.0|33|FD|1|ROIShapeControlPoints
0029|Silhouette ROI V1.0|34|UL|1|ROIDontSave
0029|Silhouette Sequence Ids V1.0|41|SQ|1|Unknown
0029|Silhouette Sequence Ids V1.0|42|SQ|1|Unknown
0029|Silhouette Sequence Ids V1.0|43|SQ|1|Unknown
0029|Silhouette V1.0|13|UL|1|Unknown
0029|Silhouette V1.0|14|UL|1|Unknown
0029|Silhouette V1.0|17|UN|1|Unknown
0029|Silhouette V1.0|18|UN|1|Unknown
0029|Silhouette V1.0|19|UL|1|Unknown
0029|Silhouette V1.0|1a|UN|1|Unknown
0029|Silhouette V1.0|1b|UL|1|Unknown
0029|Silhouette V1.0|1c|UL|1|Unknown
0029|Silhouette V1.0|1d|UN|1|Unknown
0029|Silhouette V1.0|1e|UN|1|Unknown
0029|Silhouette V1.0|21|US|1|Unknown
0029|Silhouette V1.0|22|US|1|Unknown
0029|Silhouette V1.0|23|US|1|Unknown
0029|Silhouette V1.0|24|US|1|Unknown
0029|Silhouette V1.0|25|US|1|Unknown
0029|Silhouette V1.0|27|UN|1|Unknown
0029|Silhouette V1.0|28|UN|1|Unknown
0029|Silhouette V1.0|29|UN|1|Unknown
0029|Silhouette V1.0|30|UN|1|Unknown
0029|Silhouette V1.0|52|US|1|Unknown
0029|Silhouette V1.0|53|LT|1|Unknown
0029|Silhouette V1.0|54|UN|1|Unknown
0029|Silhouette V1.0|55|LT|1|Unknown
0029|Silhouette V1.0|56|LT|1|Unknown
0029|Silhouette V1.0|57|UN|1|Unknown
0135|SONOWAND AS|10|LO|1|UltrasoundScannerName
0135|SONOWAND AS|11|LO|1|TransducerSerial
0135|SONOWAND AS|12|LO|1|ProbeApplication
0017|SVISION|00|LO|1|ExtendedBodyPart
0017|SVISION|10|LO|1|ExtendedViewPosition
0017|SVISION|F0|IS|1|ImagesSOPClass
0019|SVISION|00|IS|1|AECField
0019|SVISION|01|IS|1|AECFilmScreen
0019|SVISION|02|IS|1|AECDensity
0019|SVISION|10|IS|1|PatientThickness
0019|SVISION|18|IS|1|BeamDistance
0019|SVISION|20|IS|1|WorkstationNumber
0019|SVISION|28|IS|1|TubeNumber
0019|SVISION|30|IS|1|BuckyGrid
0019|SVISION|34|IS|1|Focus
0019|SVISION|38|IS|1|Child
0019|SVISION|40|IS|1|CollimatorDistanceX
0019|SVISION|41|IS|1|CollimatorDistanceY
0019|SVISION|50|IS|1|CentralBeamHeight
0019|SVISION|60|IS|1|BuckyAngle
0019|SVISION|68|IS|1|CArmAngle
0019|SVISION|69|IS|1|CollimatorAngle
0019|SVISION|70|IS|1|FilterNumber
0019|SVISION|74|LO|1|FilterMaterial1
0019|SVISION|75|LO|1|FilterMaterial2
0019|SVISION|A8|DS|1|ExtendedXRayTubeCurrent
0021|SVISION|00|DS|1|NoiseReduction
0021|SVISION|01|DS|1|ContrastAmplification
0021|SVISION|02|DS|1|EdgeContrastBoosting
0021|SVISION|03|DS|1|LatitudeReduction
0021|SVISION|10|LO|1|FindRangeAlgorithm
0021|SVISION|11|DS|1|ThresholdCAlgorithm
0021|SVISION|20|LO|1|SensometricCurve
0021|SVISION|30|DS|1|LowerWindowOffset
0021|SVISION|31|DS|1|UpperWindowOffset
0021|SVISION|40|DS|1|MinPrintableDensity
0021|SVISION|41|DS|1|MaxPrintableDensity
0021|SVISION|90|DS|1|Brightness
0021|SVISION|91|DS|1|Contrast
0021|SVISION|92|DS|1|ShapeFactor
0023|SVISION|00|LO|1|ImageLaterality
0023|SVISION|01|IS|1|LetterPosition
0023|SVISION|02|IS|1|BurnedInAnnotation
0023|SVISION|03|LO|1|Unknown
0023|SVISION|F0|IS|1|ImageSOPClass
0025|SVISION|00|IS|1|OriginalImage
0025|SVISION|01|IS|1|NotProcessedImage
0025|SVISION|02|IS|1|CutOutImage
0025|SVISION|03|IS|1|DuplicatedImage
0025|SVISION|04|IS|1|StoredImage
0025|SVISION|05|IS|1|RetrievedImage
0025|SVISION|06|IS|1|RemoteImage
0025|SVISION|07|IS|1|MediaStoredImage
0025|SVISION|08|IS|1|ImageState
0025|SVISION|20|LO|1|SourceImageFile
0025|SVISION|21|UI|1|Unknown
0027|SVISION|00|IS|1|NumberOfSeries
0027|SVISION|01|IS|1|NumberOfStudies
0027|SVISION|10|DT|1|OldestSeries
0027|SVISION|11|DT|1|NewestSeries
0027|SVISION|12|DT|1|OldestStudy
0027|SVISION|13|DT|1|NewestStudy
0009|TOSHIBA_MEC_1.0|01|LT|1|Unknown
0009|TOSHIBA_MEC_1.0|02|US|1-n|Unknown
0009|TOSHIBA_MEC_1.0|03|US|1-n|Unknown
0009|TOSHIBA_MEC_1.0|04|US|1-n|Unknown
0011|TOSHIBA_MEC_1.0|01|LT|1|Unknown
0011|TOSHIBA_MEC_1.0|02|US|1-n|Unknown
0019|TOSHIBA_MEC_1.0|01|US|1-n|Unknown
0019|TOSHIBA_MEC_1.0|02|US|1-n|Unknown
0021|TOSHIBA_MEC_1.0|01|US|1-n|Unknown
0021|TOSHIBA_MEC_1.0|02|US|1-n|Unknown
0021|TOSHIBA_MEC_1.0|03|US|1-n|Unknown
7ff1|TOSHIBA_MEC_1.0|01|US|1-n|Unknown
7ff1|TOSHIBA_MEC_1.0|02|US|1-n|Unknown
7ff1|TOSHIBA_MEC_1.0|03|US|1-n|Unknown
7ff1|TOSHIBA_MEC_1.0|10|US|1-n|Unknown
0019|TOSHIBA_MEC_CT_1.0|01|IS|1|Unknown
0019|TOSHIBA_MEC_CT_1.0|02|IS|1|Unknown
0019|TOSHIBA_MEC_CT_1.0|03|US|1-n|Unknown
0019|TOSHIBA_MEC_CT_1.0|04|LT|1|Unknown
0019|TOSHIBA_MEC_CT_1.0|05|LT|1|Unknown
0019|TOSHIBA_MEC_CT_1.0|06|US|1-n|Unknown
0019|TOSHIBA_MEC_CT_1.0|07|US|1-n|Unknown
0019|TOSHIBA_MEC_CT_1.0|08|LT|1|OrientationHeadFeet
0019|TOSHIBA_MEC_CT_1.0|09|LT|1|ViewDirection
0019|TOSHIBA_MEC_CT_1.0|0a|LT|1|OrientationSupineProne
0019|TOSHIBA_MEC_CT_1.0|0b|DS|1|Unknown
0019|TOSHIBA_MEC_CT_1.0|0c|US|1-n|Unknown
0019|TOSHIBA_MEC_CT_1.0|0d|TM|1|Time
0019|TOSHIBA_MEC_CT_1.0|0e|DS|1|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|01|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|02|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|03|IS|1|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|04|IS|1|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|05|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|07|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|08|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|09|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|0a|LT|1|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|0b|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|0c|US|1-n|Unknown
7ff1|TOSHIBA_MEC_CT_1.0|0d|US|1-n|Unknown
0009|ACUSON:1.2.840.113680.1.0:0910|00|IS|1|Unknown
0009|ACUSON:1.2.840.113680.1.0:0910|01|IS|1|Unknown
0009|ACUSON:1.2.840.113680.1.0:0910|02|LO|1|Patient Registration Custom Field 1
0009|ACUSON:1.2.840.113680.1.0:0910|03|LO|1|Patient Registration Custom Field 2
0009|ACUSON:1.2.840.113680.1.0:0910|04|LO|1|Indications
0009|ACUSON:1.2.840.113680.1.0:0910|0f|LT|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|02|US|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|0b|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|0c|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|20|FL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|22|FL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|00|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|01|US|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|0d|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|10|SH|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|24|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|25|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|26|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|27|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|28|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|29|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|2a|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|2b|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|2c|UL|1-n|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|30|SQ|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|31|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|32|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|33|FL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|34|FL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|35|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|36|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|37|FL|1|Unknown
0087|AGFA-AG_HPState|02|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|38|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|50|SH|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|52|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|54|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|60|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|61|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|62|FD|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|63|FD|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|64|FD|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|65|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|66|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|67|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|68|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|69|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|6a|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|6b|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|6c|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|72|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|73|FD|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|74|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|75|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|76|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|77|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|78|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|79|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7a|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7b|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7c|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7d|LO|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7e|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|7f|SL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|80|UL|1-n|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|81|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|82|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|83|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|85|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|89|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|8a|FD|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|8b|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|8c|UL|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|8d|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|86|OB|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|88|FD|1|Unknown
0087|AGFA-AG_HPState|03|SL|2|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|f1|UL|1-n|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7f10|f5|IS|1|Unknown
7fdf|ACUSON:1.2.840.113680.1.0:7ffe|00|OB|1|Unknown
0011|AgilityRuntime|20|LO|1|Unknown
0011|AgilityRuntime|21|LO|1|Unknown
0011|AgilityRuntime|22|LO|1|Unknown
0011|AGFA-AG_HPState|11|SH|1|Unknown
0019|AGFA-AG_HPState|a0|SQ|1|Unknown
0019|AGFA-AG_HPState|a1|FL|1|Unknown
0019|AGFA-AG_HPState|a2|FL|1|Unknown
0019|AGFA-AG_HPState|a3|FL|1|Unknown
0019|AGFA-AG_HPState|a4|FL|1|Unknown
0019|AGFA|05|ST|1|Cassette Data Stream
0019|AGFA|10|ST|1|Image Processing Parameters
0019|AGFA|11|LO|1|Identification Data
0019|AGFA|13|LO|1|Sensitometry Name
0019|AGFA|14|ST|1|Window Level List
0019|AGFA|15|LO|1|Dose Monitoring
0019|AGFA|16|LO|1|Other Info
0019|AGFA|1a|LO|1|Clipped Exposure Deviation
0019|AGFA|1b|LO|1|Logarithmic PLT Full Scale
0019|AGFA|60|US|1|Total Number Series
0019|AGFA|61|SH|1|Session Number
0019|AGFA|62|SH|1|ID Station Name
0019|AGFA|65|US|1|Number of Images in Study to be Transmitted
0019|AGFA|70|US|1|Total Number Images
0019|AGFA|80|ST|1|Geometrical Transformations
0019|AGFA|81|ST|1|Roam Origin
0019|AGFA|82|US|1|Zoom Factor
0019|AGFA|93|CS|1|Status
0019|AGFA_ADC_Compact|30|ST|1|Data stream from cassette
0019|AGFA_ADC_Compact|40|ST|1|Set of destination Ids
0019|AGFA_ADC_Compact|50|ST|1|Set of processing codes
0019|AGFA_ADC_Compact|60|US|1|Number of series in study
0019|AGFA_ADC_Compact|61|US|1|Session Number
0019|AGFA_ADC_Compact|62|SH|1|ID station name
0019|AGFA_ADC_Compact|70|US|1|Number of images in series
0019|AGFA_ADC_Compact|71|US|1|Break condition
0019|AGFA_ADC_Compact|72|US|1|Wait (or Hold) flag
0019|AGFA_ADC_Compact|73|US|1|ScanRes flag
0019|AGFA_ADC_Compact|74|SH|1|Operation code
0019|AGFA_ADC_Compact|95|CS|1|Image quality
0019|Agfa ADC NX|07|CS|1|Unknown
0019|Agfa ADC NX|09|SQ|1|Unknown
0019|Agfa ADC NX|21|FL|1|Unknown
0019|Agfa ADC NX|28|CS|1|Unknown
0019|Agfa ADC NX|f0|LO|1|User Defined field 1
0019|Agfa ADC NX|f1|LO|1|User Defined field 2
0019|Agfa ADC NX|f2|LO|1|User Defined field 3
0019|Agfa ADC NX|f3|LO|1|User Defined field 4
0019|Agfa ADC NX|f4|LO|1|User Defined field 5
0019|Agfa ADC NX|f5|CS|1|Cassette Orientation
0019|Agfa ADC NX|f6|DS|1|Plate Sensitivity
0019|Agfa ADC NX|f7|DS|1|Plate Erasability
0019|Agfa ADC NX|f8|IS|1|Unknown
0019|Agfa ADC NX|fa|IS|1|Unknown
0019|Agfa ADC NX|fc|IS|1|Unknown
0019|Agfa ADC NX|fd|CS|1|Unknown
0019|Agfa ADC NX|fe|CS|1|Unknown
0031|AGFA PACS Archive Mirroring 1.0|00|CS|1|Unknown
0031|AGFA PACS Archive Mirroring 1.0|01|UL|1|Unknown
0029|MITRA PRESENTATION 1.0|00|CS|1|Rotation
0029|MITRA PRESENTATION 1.0|01|LO|1|Window Width
0029|MITRA PRESENTATION 1.0|02|LO|1|Window Centre
0029|MITRA PRESENTATION 1.0|03|IS|1|Invert
0029|MITRA PRESENTATION 1.0|04|IS|1|Has Tabstop
0029|MITRA PRESENTATION 1.0|05|CS|1|Smooth Rotation
0029|MITRA PRESENTATION 1.0|10|CS|1|Unknown
0029|MITRA PRESENTATION 1.0|11|CS|1|Unknown
0029|MITRA PRESENTATION 1.0|12|CS|1|Unknown
0029|MITRA PRESENTATION 1.0|13|CS|1|Unknown
0029|MITRA OBJECT DOCUMENT 1.0|00|OB|1|IMPAX Object Document
0029|MITRA OBJECT DOCUMENT 1.0|01|OB|1|IMPAX Markup XML Stored
0029|MITRA MARKUP 1.0|00|OB|1-n|Markup1
0029|MITRA MARKUP 1.0|01|OB|1-n|Markup2
0029|MITRA MARKUP 1.0|02|OB|1-n|Markup3
0029|MITRA MARKUP 1.0|03|OB|1-n|Markup4
0029|MITRA MARKUP 1.0|04|OB|1-n|Markup5
0029|MITRA MARKUP 1.0|05|OB|1-n|Markup6
0029|MITRA MARKUP 1.0|06|OB|1-n|Markup7
0029|MITRA MARKUP 1.0|07|OB|1-n|Markup8
0029|MITRA MARKUP 1.0|08|OB|1-n|Markup9
0029|MITRA MARKUP 1.0|09|OB|1-n|Markup10
0029|MITRA MARKUP 1.0|10|OB|1-n|Markup11
0029|MITRA MARKUP 1.0|11|OB|1-n|Markup12
0029|MITRA MARKUP 1.0|12|OB|1-n|Markup13
0029|MITRA MARKUP 1.0|13|OB|1-n|Markup14
0029|MITRA MARKUP 1.0|14|OB|1-n|Markup14
0029|AgilityRuntime|11|CS|1|Unknown
0029|AgilityRuntime|12|US|1|Unknown
0029|AgilityRuntime|13|US|1|Unknown
0029|AgilityRuntime|14|US|1|Unknown
0029|AgilityRuntime|1f|US|1|Unknown
0031|MITRA LINKED ATTRIBUTES 1.0|20|IS|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|02|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|04|CS|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|06|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|08|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|0a|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|0c|LO|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|0e|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|13|PN|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|14|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|15|OB|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|16|PN|1|Unknown
0033|MITRA OBJECT UTF8 ATTRIBUTES 1.0|19|PN|1|Unknown
0033|MITRA OBJECT ATTRIBUTES 1.0|02|LO|1|Unknown
0033|MITRA OBJECT ATTRIBUTES 1.0|04|LO|1|Unknown
0033|MITRA OBJECT ATTRIBUTES 1.0|06|LO|1|Unknown
0033|MITRA OBJECT ATTRIBUTES 1.0|08|LO|1|Unknown
0087|AGFA-AG_HPState|04|SL|2|Unknown
0033|MITRA OBJECT ATTRIBUTES 1.0|0a|LO|1|Unknown
0071|AGFA-AG_HPState|18|SQ|1|Unknown
0071|AGFA-AG_HPState|19|SQ|1|Unknown
0071|AGFA-AG_HPState|1a|SQ|1|Unknown
0071|AGFA-AG_HPState|1c|SQ|1|Unknown
0071|AGFA-AG_HPState|1e|SQ|1|Unknown
0071|AGFA-AG_HPState|20|FL|1-n|Unknown
0071|AGFA-AG_HPState|21|FD|1-n|Unknown
0071|AGFA-AG_HPState|22|FD|1-n|Unknown
0071|AGFA-AG_HPState|23|FD|1-n|Unknown
0071|AGFA-AG_HPState|24|FD|1|Unknown
0071|AGFA-AG_HPState|2b|FD|1-n|Unknown
0071|AGFA-AG_HPState|2c|FD|3|Unknown
0071|AGFA-AG_HPState|2d|FD|1|Unknown
0071|AgilityOverlay|01|ST|1|Unknown
0071|AgilityOverlay|02|ST|1|Unknown
0071|AgilityOverlay|03|ST|1|Unknown
0071|AgilityOverlay|05|ST|1|Unknown
0071|AgilityOverlay|06|SQ|1|Unknown
0071|AgilityOverlay|07|ST|1|Unknown
0071|AgilityOverlay|08|CS|1|Unknown
0071|AgilityOverlay|09|ST|1|Unknown
0071|AgilityOverlay|0a|CS|1|Unknown
0071|AgilityOverlay|10|FL|1|Unknown
0071|AgilityOverlay|11|ST|1|Unknown
0071|AgilityOverlay|12|CS|1|Unknown
0071|AgilityOverlay|13|US|1|Unknown
0071|AgilityOverlay|14|US|1|Unknown
0071|AgilityOverlay|15|FD|1-n|Unknown
0071|AgilityOverlay|16|ST|1|Unknown
0071|AgilityOverlay|17|ST|1|Unknown
0071|AgilityOverlay|18|CS|1|Unknown
0071|AgilityOverlay|19|ST|1|Unknown
0071|AgilityOverlay|1b|ST|1|Unknown
0071|AgilityOverlay|1c|ST|1|Unknown
0071|AgilityOverlay|1d|ST|1|Unknown
0071|AgilityOverlay|22|ST|1|Unknown
0071|AgilityOverlay|2c|ST|1|Unknown
0071|AgilityOverlay|2d|SQ|1|Unknown
0071|AgilityOverlay|2e|US|1|Unknown
0071|AgilityOverlay|50|CS|1|Unknown
0071|AgilityOverlay|51|CS|1|Unknown
0071|AgilityOverlay|52|LT|1|Unknown
0071|AgilityOverlay|53|CS|1|Unknown
0071|AgilityOverlay|54|CS|1|Unknown
0071|AgilityOverlay|55|CS|1|Unknown
0071|AgilityOverlay|56|CS|1|Unknown
0071|AgilityOverlay|57|CS|1|Unknown
0071|AgilityOverlay|59|FL|1|Unknown
0071|AgilityOverlay|5a|FL|1|Unknown
0071|AgilityOverlay|5b|FL|2|Unknown
0071|AgilityOverlay|5c|FL|4|Unknown
0071|AgilityOverlay|5d|CS|1|Unknown
0071|AgilityOverlay|60|FD|1|Unknown
0073|AGFA-AG_HPState|23|SH|1|Unknown
0073|AGFA-AG_HPState|24|SQ|1|Unknown
0073|AGFA-AG_HPState|28|SQ|1|Unknown
0073|AGFA-AG_HPState|80|FL|1|Unknown
0075|AGFA-AG_HPState|10|LO|1|Unknown
0087|AGFA-AG_HPState|01|LO|1|Unknown
0087|AGFA-AG_HPState|05|FD|2|Unknown
0087|AGFA-AG_HPState|06|FD|2|Unknown
0087|AGFA-AG_HPState|07|FD|2|Unknown
0087|AGFA-AG_HPState|08|FD|2|Unknown
0035|AGFA KOSD 1.0|00|SH|1|Unknown
0035|AGFA KOSD 1.0|03|LT|1|Unknown
2e13|agfa/displayableImages|10|IS|1|Unknown
2e13|agfa/displayableImages|11|IS|1|Unknown
7fdb|agfa/xeroverse|99|LO|1|Unknown
0009|Camtronics image level data|04|IS|1|Unknown
0009|Camtronics image level data|06|IS|1|Unknown
0009|Camtronics image level data|09|LO|1|Unknown
0009|Camtronics image level data|16|AE|1|Unknown
0009|Camtronics image level data|17|CS|1|Unknown
0009|Camtronics image level data|18|IS|1|Unknown
0009|QCA Results|00|CS|1|Analysis Type
0009|QCA Results|04|LO|1|Segment Name
0009|QCA Results|12|DS|1|Pre-procedure Catheter Size
0009|QCA Results|13|DS|1|Pre-procedure Reference Diameter
0009|QCA Results|14|DS|1|Pre-procedure Minimum Lumen Diameter
0009|QCA Results|15|DS|1|Pre-procedure Average Diameter
0009|QCA Results|16|DS|1|Pre-procedure Stenosis Length
0009|QCA Results|17|DS|1|Pre-procedure Stenosis %
0009|QCA Results|18|DS|1|Pre-procedure Geometric Area Reduction %
0009|QCA Results|22|DS|1|Post-procedure Catheter Size
0009|QCA Results|23|DS|1|Post-procedure Reference Diameter
0009|QCA Results|24|DS|1|Post-procedure Minimum Lumen Diameter
0009|QCA Results|25|DS|1|Post-procedure Average Diameter
0009|QCA Results|26|DS|1|Post-procedure Stenosis Length
0009|QCA Results|27|DS|1|Post-procedure Stenosis %
0009|QCA Results|28|DS|1|Post-procedure Geometric Area Reduction %
0003|ELSCINT1|01|OW|1|Offset List Structure
00e1|ELSCINT1|01|US|1|Data Dictionary Version
00e1|ELSCINT1|05|IS|1|Unknown
00e1|ELSCINT1|06|IS|1|Unknown
00e1|ELSCINT1|07|IS|1|Unknown
00e1|ELSCINT1|14|CS|1|Unknown
00e1|ELSCINT1|18|OB|1|Unknown
0119|MRSC|11a1|IS|1|PhantCalibNParms
00e1|ELSCINT1|22|DS|2|Presentation Relative Center
00e1|ELSCINT1|23|DS|2|Presentation Relative Part
00e1|ELSCINT1|24|CS|1|Unknown
00e1|ELSCINT1|25|CS|1|Unknown
00e1|ELSCINT1|30|UI|1|Unknown
00e1|ELSCINT1|31|CS|1|Unknown
00e1|ELSCINT1|32|US|2|Unknown
00e1|ELSCINT1|37|DS|1|Total Dose Savings
00e1|ELSCINT1|39|SQ|1|Unknown
00e1|ELSCINT1|3e|IS|1|Unknown
00e1|ELSCINT1|3f|CS|1|Unknown
00e1|ELSCINT1|40|SH|1|Image Label
00e1|ELSCINT1|41|DS|1|Unknown
00e1|ELSCINT1|42|LO|1|Unknown
00e1|ELSCINT1|43|IS|1|Unknown
00e1|ELSCINT1|50|DS|1|Acquisition Duration
00e1|ELSCINT1|51|SH|1|Unknown
00e1|ELSCINT1|60|CS|1|Unknown
00e1|ELSCINT1|61|LO|1|Protocol File Name
00e1|ELSCINT1|62|CS|1|Unknown
00e1|ELSCINT1|63|SH|1|Patient Language
00e1|ELSCINT1|65|LO|1|Unknown
00e1|ELSCINT1|6a|IS|1|Unknown
00e1|ELSCINT1|6b|IS|1|Unknown
00e1|ELSCINT1|a0|LO|1|Unknown
00e1|ELSCINT1|c4|DS|1|Unknown
00e1|ELSCINT1|cf|IS|1|Unknown
00e1|ELSCINT1|eb|US|1|Unknown
00e1|ELSCINT1|ec|US|1|Unknown
01e1|ELSCINT1|18|OB|1|Unknown
01e1|ELSCINT1|21|ST|1|Unknown
01e1|ELSCINT1|26|CS|1|Phantom Type
01e1|ELSCINT1|34|IS|1|Unknown
01e1|ELSCINT1|40|UI|1|Unknown
01e1|ELSCINT1|41|OW|1|Unknown
01f1|ELSCINT1|01|CS|1|Acquisition Type
01f1|ELSCINT1|02|CS|1|Focal Spot Resolution
01f1|ELSCINT1|03|CS|1|Concurrent Slices Generation
01f1|ELSCINT1|04|CS|1|Angular Sampling Density
01f1|ELSCINT1|05|DS|1|Reconstruction Arc
01f1|ELSCINT1|07|DS|1|Table Velocity
01f1|ELSCINT1|08|DS|1|Acquisition Length
01f1|ELSCINT1|0a|US|1|Edge Enhancement Weight
01f1|ELSCINT1|0c|DS|1|Scanner Relative Center
01f1|ELSCINT1|0d|DS|1|Rotation Angle
01f1|ELSCINT1|0e|FL|1|Unknown
01f1|ELSCINT1|26|DS|1|Pitch
01f1|ELSCINT1|27|DS|1|Rotation Time
01f1|ELSCINT1|28|DS|1|Table Increment
01f1|ELSCINT1|30|US|1|Unknown
01f1|ELSCINT1|32|CS|1|Image View Convention
01f1|ELSCINT1|33|DS|1|Cycle Time
01f1|ELSCINT1|36|CS|1|Unknown
01f1|ELSCINT1|37|DS|1|Unknown
01f1|ELSCINT1|38|LO|1|Unknown
01f1|ELSCINT1|39|LO|1|Unknown
01f1|ELSCINT1|40|CS|1|Unknown
01f1|ELSCINT1|42|SH|1|Unknown
01f1|ELSCINT1|43|LO|1|Unknown
01f1|ELSCINT1|44|OW|1|Unknown
01f1|ELSCINT1|45|IS|1|Unknown
01f1|ELSCINT1|46|FL|1|Unknown
01f1|ELSCINT1|47|SH|1|Unknown
01f1|ELSCINT1|49|DS|1|Unknown
01f1|ELSCINT1|4a|SH|1|Unknown
01f1|ELSCINT1|4b|SH|1|Unknown
01f1|ELSCINT1|4c|SH|1|Unknown
01f1|ELSCINT1|4d|SH|1|Unknown
01f1|ELSCINT1|4e|LO|1|Unknown
01f1|ELSCINT1|53|SH|1|Unknown
01f3|ELSCINT1|01|SQ|1|Unknown
01f3|ELSCINT1|02|SS|1|Unknown
01f3|ELSCINT1|03|FL|2|Unknown
01f3|ELSCINT1|04|FL|1|Unknown
01f3|ELSCINT1|11|SQ|1|Unknown
01f3|ELSCINT1|12|SS|1|Unknown
01f3|ELSCINT1|13|FL|2|Unknown
01f3|ELSCINT1|14|FL|1|Unknown
01f3|ELSCINT1|15|US|1|Unknown
01f3|ELSCINT1|16|FL|1|Unknown
01f3|ELSCINT1|17|FL|1|Unknown
01f3|ELSCINT1|18|SH|1|Unknown
01f3|ELSCINT1|19|FL|1|Unknown
01f3|ELSCINT1|23|US|1|Unknown
01f3|ELSCINT1|24|IS|2|Unknown
01f7|ELSCINT1|10|OB|1|Unknown
01f7|ELSCINT1|11|OW|1|Unknown
01f7|ELSCINT1|13|OW|1|Unknown
01f7|ELSCINT1|14|OW|1|Unknown
01f7|ELSCINT1|15|OW|1|Unknown
01f7|ELSCINT1|16|OW|1|Unknown
01f7|ELSCINT1|17|OW|1|Unknown
01f7|ELSCINT1|18|OW|1|Unknown
01f7|ELSCINT1|19|OW|1|Unknown
01f7|ELSCINT1|1a|OW|1|Unknown
01f7|ELSCINT1|1b|OW|1|Unknown
01f7|ELSCINT1|1c|OW|1|Unknown
01f7|ELSCINT1|1e|OW|1|Unknown
01f7|ELSCINT1|1f|OW|1|Unknown
01f7|ELSCINT1|22|UI|1|Unknown
01f7|ELSCINT1|23|OW|1|Unknown
01f7|ELSCINT1|25|OW|1|Unknown
01f7|ELSCINT1|26|OW|1|Unknown
01f7|ELSCINT1|27|OW|1|Unknown
01f7|ELSCINT1|28|OW|1|Unknown
01f7|ELSCINT1|29|OW|1|Unknown
01f7|ELSCINT1|2b|OW|1|Unknown
01f7|ELSCINT1|2c|OW|1|Unknown
01f7|ELSCINT1|2d|OW|1|Unknown
01f7|ELSCINT1|2e|OW|1|Unknown
01f7|ELSCINT1|30|OW|1|Unknown
01f7|ELSCINT1|31|OW|1|Unknown
01f7|ELSCINT1|5c|OW|1|Unknown
01f7|ELSCINT1|70|OW|1|Unknown
01f7|ELSCINT1|73|OW|1|Unknown
01f7|ELSCINT1|74|OW|1|Unknown
01f7|ELSCINT1|75|OW|1|Unknown
01f7|ELSCINT1|7f|OW|1|Unknown
01f9|ELSCINT1|01|LO|1|SP Filter
01f9|ELSCINT1|04|IS|1|Adaptive Filter
01f9|ELSCINT1|05|IS|1|Recon Increment
01f9|ELSCINT1|08|DS|1|Unknown
01f9|ELSCINT1|09|DS|1|Unknown
07a1|ELSCINT1|02|UL|1|Unknown
07a1|ELSCINT1|07|US|3|Unknown
07a1|ELSCINT1|08|DS|1-n|Unknown
07a1|ELSCINT1|09|OW|1|Unknown
07a1|ELSCINT1|0a|OB|1|Unknown
07a1|ELSCINT1|0c|US|1|Unknown
07a1|ELSCINT1|10|LO|1|Unknown
07a1|ELSCINT1|11|CS|1|Unknown
07a1|ELSCINT1|12|FL|1-n|Unknown
07a1|ELSCINT1|13|UL|1|Unknown
07a1|ELSCINT1|16|FL|1-n|Unknown
07a1|ELSCINT1|18|SQ|1|Unknown
07a1|ELSCINT1|19|FL|1|Unknown
07a1|ELSCINT1|1c|FL|1-n|Unknown
07a1|ELSCINT1|2a|CS|1|Unknown
07a1|ELSCINT1|2b|CS|1|Unknown
07a1|ELSCINT1|36|AE|1|Unknown
07a1|ELSCINT1|3d|US|1|Unknown
07a1|ELSCINT1|40|CS|1|Unknown
07a1|ELSCINT1|43|IS|1|Unknown
07a1|ELSCINT1|47|CS|1|Unknown
07a1|ELSCINT1|50|US|1|Unknown
07a1|ELSCINT1|56|US|1|Unknown
07a1|ELSCINT1|70|SH|1|Unknown
07a1|ELSCINT1|71|SH|1|Unknown
07a1|ELSCINT1|75|LO|2|Unknown
07a1|ELSCINT1|85|UL|1|Unknown
07a1|ELSCINT1|87|LT|1|Unknown
07a1|ELSCINT1|88|CS|1|Unknown
07a1|ELSCINT1|98|CS|1|Unknown
07a1|ELSCINT1|9f|CS|1|Unknown
07a3|ELSCINT1|01|LO|1|Unknown
07a3|ELSCINT1|03|CS|1|Unknown
07a3|ELSCINT1|05|CS|1|Unknown
07a3|ELSCINT1|06|CS|1|Unknown
07a3|ELSCINT1|13|SH|1|Unknown
07a3|ELSCINT1|14|ST|1|Unknown
07a3|ELSCINT1|15|ST|1|Unknown
07a3|ELSCINT1|17|SH|1|Unknown
07a3|ELSCINT1|1b|ST|1|Unknown
07a3|ELSCINT1|1f|ST|1|Unknown
07a3|ELSCINT1|22|ST|1|Unknown
07a3|ELSCINT1|23|ST|1|Unknown
07a3|ELSCINT1|34|SH|1|Unknown
07a3|ELSCINT1|43|DS|1-n|Unknown
07a3|ELSCINT1|55|SH|1|Unknown
07a3|ELSCINT1|61|LT|1|Unknown
07a3|ELSCINT1|62|SQ|1|Unknown
07a3|ELSCINT1|63|SQ|1|Unknown
07a3|ELSCINT1|64|IS|1-n|Unknown
07a3|ELSCINT1|65|CS|1|Unknown
07a3|ELSCINT1|66|IS|1|Unknown
07a3|ELSCINT1|80|SQ|1|Unknown
07a3|ELSCINT1|99|CS|1|Unknown
07a3|ELSCINT1|9c|CS|1|Unknown
07a3|ELSCINT1|9f|CS|1|Unknown
07a3|ELSCINT1|b9|CS|1|Unknown
07a3|ELSCINT1|bb|CS|1|Unknown
07a5|ELSCINT1|00|LO|1|Unknown
07a5|ELSCINT1|56|CS|1|Unknown
5001|ELSCINT1|70|SQ|1|Unknown
5001|ELSCINT1|71|SH|1|Unknown
5001|ELSCINT1|80|SQ|1|Unknown
5001|ELSCINT1|81|SH|1|Unknown
5001|ELSCINT1|82|US|3|Unknown
5001|ELSCINT1|83|FL|1-n|Unknown
5001|ELSCINT1|84|SQ|1|Unknown
7fdf|ELSCINT1|f0|OB|1|Unknown
7fdf|ELSCINT1|ff|SH|1|Unknown
0009|GEMS_PETD_01|02|LO|1|Patient ID
0009|GEMS_PETD_01|03|SH|1|Patient Compatible Version
0009|GEMS_PETD_01|04|SH|1|Patient Software Version
0009|GEMS_PETD_01|05|DT|1|Patient DateTime
0009|GEMS_PETD_01|06|SL|1|Patient Type
0009|GEMS_PETD_01|07|UI|1|Exam ID
0009|GEMS_PETD_01|08|SH|1|Exam Compatible Version
0009|GEMS_PETD_01|09|SH|1|Exam Software Version
0009|GEMS_PETD_01|0a|UI|1|Scan ID
0009|GEMS_PETD_01|0c|SH|1|Scan Software Version
0009|GEMS_PETD_01|0d|DT|1|Scan Date Time
0009|GEMS_PETD_01|0e|DT|1|Scan Ready
0009|GEMS_PETD_01|0f|ST|1|Scan Description
0009|GEMS_PETD_01|10|LO|1|Hospital Name
0009|GEMS_PETD_01|11|LO|1|Scanner Description
0009|GEMS_PETD_01|12|LO|1|Manufacturer
0009|GEMS_PETD_01|13|UI|1|FOR Identifier
0009|GEMS_PETD_01|14|LO|1|Landmark Name
0009|GEMS_PETD_01|15|SH|1|Landmark Abbrev
0009|GEMS_PETD_01|16|SL|1|Patient Position
0009|GEMS_PETD_01|17|SL|1|Scan Perspective
0009|GEMS_PETD_01|18|SL|1|Scan Type
0009|GEMS_PETD_01|19|SL|1|Scan Mode
0009|GEMS_PETD_01|1a|SL|1|Start Condition
0009|GEMS_PETD_01|1b|SL|1|Start Condition Data
0009|GEMS_PETD_01|1c|SL|1|Sel Stop Condition
0009|GEMS_PETD_01|1d|SL|1|Sel Stop Condition Data
0009|GEMS_PETD_01|1e|SL|1|Collect Deadtime
0009|GEMS_PETD_01|1f|SL|1|Collect Singles
0009|GEMS_PETD_01|20|SL|1|Collect Count Rate
0119|MRSC|11a2|DS|1-n|PhantCalibParam
0009|GEMS_PETD_01|22|SL|1|Delayed Events
0009|GEMS_PETD_01|23|SL|1|Delayed Bias
0009|GEMS_PETD_01|24|SL|1|Word Size
0009|GEMS_PETD_01|25|SL|1|Axial Acceptance
0009|GEMS_PETD_01|26|SL|1|Axial Angle 3D
0009|GEMS_PETD_01|27|SL|1|Theta Compression
0009|GEMS_PETD_01|28|SL|1|Axial Compression
0009|GEMS_PETD_01|2a|SL|1|Collimation
0009|GEMS_PETD_01|2b|SL|1|Scan FOV
0009|GEMS_PETD_01|2c|SL|1|Axial FOV
0009|GEMS_PETD_01|2d|SL|1|Event Separation
0009|GEMS_PETD_01|2e|SL|1|Mask Width
0009|GEMS_PETD_01|2f|SL|1|Binning Mode
0009|GEMS_PETD_01|30|SL|1|Trig Rej Method
0009|GEMS_PETD_01|31|SL|1|Number For Reject
0009|GEMS_PETD_01|32|SL|1|Lower Reject Limit
0009|GEMS_PETD_01|33|SL|1|Upper Reject Limit
0009|GEMS_PETD_01|34|SL|1|Triggers Acquired
0009|GEMS_PETD_01|35|SL|1|Triggers Rejected
0009|GEMS_PETD_01|36|LO|1|Tracer Name
0009|GEMS_PETD_01|37|LO|1|Batch Description
0009|GEMS_PETD_01|38|FL|1|Tracer Activity
0009|GEMS_PETD_01|39|DT|1|Measured Date Time
0009|GEMS_PETD_01|3a|FL|1|Pre Inj Volume
0009|GEMS_PETD_01|3b|DT|1|Administered Date Time
0009|GEMS_PETD_01|3d|DT|1|Post Injected Date Time
0009|GEMS_PETD_01|3e|SH|1|Radio Nuclide Name
0009|GEMS_PETD_01|3f|FL|1|Half Life
0009|GEMS_PETD_01|40|FL|1|Positron Fraction
0009|GEMS_PETD_01|41|SL|1|Source 1 Holder
0009|GEMS_PETD_01|42|FL|1|Source 1 Activity
0009|GEMS_PETD_01|43|DT|1|Source 1 Meas DT
0009|GEMS_PETD_01|44|SH|1|Source 1 Radio Nuclide
0009|GEMS_PETD_01|45|FL|1|Source 1 Half Life
0009|GEMS_PETD_01|46|SL|1|Source 2 Holder
0009|GEMS_PETD_01|47|FL|1|Source 2 Activity
0009|GEMS_PETD_01|48|DT|1|Source 2 Meas DT
0009|GEMS_PETD_01|49|SH|1|Source 2 Radio Nuclide
0009|GEMS_PETD_01|4a|FL|1|Source 2 Half Life
0009|GEMS_PETD_01|4b|SL|1|Source Speed
0009|GEMS_PETD_01|4c|FL|1|Source Location
0009|GEMS_PETD_01|4d|SL|1|Emission Present
0009|GEMS_PETD_01|4e|SL|1|Lower Axial Acc
0009|GEMS_PETD_01|4f|SL|1|Upper Axial Acc
0009|GEMS_PETD_01|50|SL|1|Lower Coinc Limit
0009|GEMS_PETD_01|52|SL|1|Coinc Delay Offset
0009|GEMS_PETD_01|53|SL|1|Coinc Output Mode
0009|GEMS_PETD_01|54|SL|1|Upper Energy Limit
0009|GEMS_PETD_01|55|SL|1|Lower Energy Limit
0009|GEMS_PETD_01|56|UI|1|Normal Cal ID
0009|GEMS_PETD_01|57|UI|1|Normal 2D Cal ID
0009|GEMS_PETD_01|58|UI|1|Blank Cal ID
0009|GEMS_PETD_01|59|UI|1|WC Cal ID
0009|GEMS_PETD_01|5a|SL|1|Derived
0009|GEMS_PETD_01|5b|LO|1|Contrast Agent
0009|GEMS_PETD_01|5c|UI|1|frame_id
0009|GEMS_PETD_01|5d|UI|1|scan_id
0119|MRSC|11a3|IS|1-n|PhantGoodFlags
0009|GEMS_PETD_01|5f|LO|1|patient_id
0009|GEMS_PETD_01|61|SH|1|software_version
0009|GEMS_PETD_01|62|ST|1|where_is_frame
0009|GEMS_PETD_01|63|SL|1|frame_size
0009|GEMS_PETD_01|64|SL|1|file_exists
0009|GEMS_PETD_01|65|SL|1|patient_entry
0009|GEMS_PETD_01|66|FL|1|table_height
0009|GEMS_PETD_01|67|FL|1|table_z_position
0009|GEMS_PETD_01|68|DT|1|landmark_datetime
0009|GEMS_PETD_01|69|SL|1|slice_count
0009|GEMS_PETD_01|6a|FL|1|start_location
0009|GEMS_PETD_01|6b|SL|1|acq_delay
0009|GEMS_PETD_01|6c|DT|1|acq_start
0009|GEMS_PETD_01|6d|SL|1|acq_duration
0009|GEMS_PETD_01|6e|SL|1|acq_bin_dur
0009|GEMS_PETD_01|6f|SL|1|acq_bin_start
0009|GEMS_PETD_01|70|SL|1|actual_stop_cond
0009|GEMS_PETD_01|71|FD|1|total_prompts
0009|GEMS_PETD_01|72|FD|1|total_delays
0009|GEMS_PETD_01|73|SL|1|frame_valid
0009|GEMS_PETD_01|74|SL|1|validity_info
0009|GEMS_PETD_01|75|SL|1|archived
0009|GEMS_PETD_01|76|SL|1|compression
0009|GEMS_PETD_01|77|SL|1|uncompressed_size
0009|GEMS_PETD_01|78|SL|1|accum_bin_dur
0009|GEMS_PETD_01|7a|SH|1|Image Set Software Version
0009|GEMS_PETD_01|7b|DT|1|Image Set Date Time
0009|GEMS_PETD_01|7c|SL|1|Image Set Source
0009|GEMS_PETD_01|7d|SL|1|Image Set Contents
0009|GEMS_PETD_01|7e|SL|1|Image Set Type
0009|GEMS_PETD_01|7f|DS|1|Image Set Reference
0009|GEMS_PETD_01|80|SL|1|Multi Patient
0009|GEMS_PETD_01|81|SL|1|Number of Normals
0009|GEMS_PETD_01|82|UI|1|Color Map ID
0009|GEMS_PETD_01|83|SL|1|Window Level Type
0009|GEMS_PETD_01|84|FL|1|Rotate
0009|GEMS_PETD_01|85|SL|1|Flip
0009|GEMS_PETD_01|86|FL|1|Zoom
0009|GEMS_PETD_01|87|SL|1|PanX
0009|GEMS_PETD_01|88|SL|1|PanY
0009|GEMS_PETD_01|89|FL|1|Window Level Min
0009|GEMS_PETD_01|8a|FL|1|Window Level Max
0009|GEMS_PETD_01|8b|SL|1|ReconMethod
0009|GEMS_PETD_01|8c|SL|1|Attenuation
0009|GEMS_PETD_01|8d|FL|1|Attenuation Coefficient
0009|GEMS_PETD_01|8e|SL|1|BP Filter
0009|GEMS_PETD_01|8f|FL|1|BP Filter Cutoff
0009|GEMS_PETD_01|90|SL|1|BP Filter Order
0009|GEMS_PETD_01|91|FL|1|BP Filter Center I
0009|GEMS_PETD_01|92|FL|1|BP Filter Center P
0009|GEMS_PETD_01|93|SL|1|Atten Smooth
0009|GEMS_PETD_01|95|SL|1|Angle Smooth Param
0009|GEMS_PETD_01|96|UI|1|Well CounterCal ID
0009|GEMS_PETD_01|97|UI|1|Trans Scan ID
0009|GEMS_PETD_01|98|UI|1|Norm Cal ID
0009|GEMS_PETD_01|99|UI|1|Blnk Cal ID
0009|GEMS_PETD_01|9a|FL|1|CAC Edge Threshold
0009|GEMS_PETD_01|9c|UI|1|Emiss Sub ID
0009|GEMS_PETD_01|9d|SS|1|Radial Filter 3D
0009|GEMS_PETD_01|9e|FL|1|Radial Cutoff 3D
0009|GEMS_PETD_01|a0|FL|1|Axial Cutoff 3D
0009|GEMS_PETD_01|a1|FL|1|Axial Start
0009|GEMS_PETD_01|a2|FL|1|Axial Spacing
0009|GEMS_PETD_01|a3|SL|1|Axial Angles Used
0009|GEMS_PETD_01|a4|SH|1|compatible_version
0009|GEMS_PETD_01|a5|SH|1|software_version
0009|GEMS_PETD_01|a6|SL|1|slice_number
0009|GEMS_PETD_01|a7|FL|1|total_counts
0009|GEMS_PETD_01|a8|OB|1|other_atts
0009|GEMS_PETD_01|a9|SL|1|other_atts_size
0009|GEMS_PETD_01|aa|SL|1|archived
0009|GEMS_PETD_01|ab|FL|1|bp_center_x
0009|GEMS_PETD_01|ac|FL|1|bp_center_y
0009|GEMS_PETD_01|ad|UI|1|trans_frame_id
0009|GEMS_PETD_01|ae|UI|1|tpluse_frame_id
0009|GEMS_PETD_01|b1|FL|1|profile_spacing
0009|GEMS_PETD_01|b2|SS|1|IR Num Iterations
0009|GEMS_PETD_01|b3|SS|1|IR Num Subsets
0009|GEMS_PETD_01|b4|FL|1|IR Recon FOV
0009|GEMS_PETD_01|b5|SS|1|IR Corr Model
0009|GEMS_PETD_01|b7|FL|1|IR Pre Filt Param
0009|GEMS_PETD_01|b8|FL|1|IR Loop Filt Param
0009|GEMS_PETD_01|b9|FL|1|Response Filt Param
0009|GEMS_PETD_01|ba|SS|1|Post Filter
0009|GEMS_PETD_01|bb|FL|1|Post Filter Param
0009|GEMS_PETD_01|bc|SS|1|IR Regularize
0009|GEMS_PETD_01|bd|FL|1|IR Regularize Param
0009|GEMS_PETD_01|be|SS|1|AC BP Filter
0009|GEMS_PETD_01|bf|FL|1|AC BP Filt Cutoff
0009|GEMS_PETD_01|c0|SL|1|AC BP Filt Order
0009|GEMS_PETD_01|c1|SS|1|AC Img Smooth
0009|GEMS_PETD_01|c2|FL|1|AC Img Smooth Parm
0009|GEMS_PETD_01|c3|SL|1|Scatter Method
0009|GEMS_PETD_01|c4|SS|1|Scatter Num Iter
0009|GEMS_PETD_01|c5|FL|1|Scatter Parm
0009|GEMS_PETD_01|c6|FL|1|seg_qc_parm
0009|GEMS_PETD_01|c7|SL|1|overlap
0009|GEMS_PETD_01|c8|UI|1|ovlp_frm_id
0009|GEMS_PETD_01|c9|UI|1|ovlp_trans_frm_id
0009|GEMS_PETD_01|ca|UI|1|ovlp_tpulse_frm_id
0009|GEMS_PETD_01|cb|FL|1|vqc_x_axis_trans
0009|GEMS_PETD_01|cc|FL|1|vqc_x_axis_tilt
0009|GEMS_PETD_01|ce|FL|1|vqc_y_axis_swivel
0009|GEMS_PETD_01|cf|FL|1|vqc_z_axis_trans
0009|GEMS_PETD_01|d0|FL|1|vqc_z_axis_roll
0009|GEMS_PETD_01|d1|LO|1|ctac_conv_scale
0009|GEMS_PETD_01|d2|UI|1|image_set_id
0009|GEMS_PETD_01|d3|SL|1|contrast_route
0009|GEMS_PETD_01|d4|LO|1|ctac_conv_scale
0009|GEMS_PETD_01|d5|FL|1|loop_filter_parm
0009|GEMS_PETD_01|d6|FL|1|image_one_loc
0009|GEMS_PETD_01|d7|FL|1|image_index_loc
0009|GEMS_PETD_01|d8|SL|1|frame_number
0009|GEMS_PETD_01|d9|SL|1|list_file_exists
0119|MRSC|11a4|DS|1-n|PhantValues
0011|GEMS_PETD_01|18|OB|1|Unknown
0023|GEMS_PETD_01|01|OB|1|raw_data_blob
5001|GEMS_PETD_01|01|UI|1|Curve ID
0009|GEMS_PETD_01|dc|FL|1|ir_z_filter_ratio
0009|GEMS_PETD_01|dd|US|1|num_of_rr_interval
0009|GEMS_PETD_01|de|US|1|num_of_time_slots
0009|GEMS_PETD_01|df|US|1|num_of_slices
0009|GEMS_PETD_01|e0|US|1|num_of_time_slices
0009|GEMS_PETD_01|e1|SL|1|unlisted_scan
0009|GEMS_PETD_01|e2|SL|1|rest_stress
0009|GEMS_PETD_01|e3|FL|1|phase percentage
0009|GEMS_PETD_01|e4|ST|1|Unknown
0009|GEMS_PETD_01|e5|FL|1|left shift
0009|GEMS_PETD_01|e6|FL|1|posterior shift
0009|GEMS_PETD_01|e7|FL|1|superior shift
0009|GEMS_PETD_01|e8|SL|1|acq_bin_num
0009|GEMS_PETD_01|e9|FL|1|acq_bin_dur_percent
0009|GEMS_PETD_01|ea|SL|1|Unknown
0009|GEMS_PETD_01|eb|FL|1|Unknown
0009|GEMS_PETD_01|ec|SL|1|Unknown
0011|GEMS_PETD_01|01|SQ|1|Unknown
0013|GEMS_PETD_01|01|SQ|1|Unknown
0017|GEMS_PETD_01|01|UI|1|correction_cal_id
0017|GEMS_PETD_01|03|SH|1|software_version
0017|GEMS_PETD_01|04|DT|1|cal_datetime
0017|GEMS_PETD_01|05|LO|1|cal_datetime
0017|GEMS_PETD_01|06|SL|1|cal_type
0017|GEMS_PETD_01|07|ST|1|where_is_corr
0017|GEMS_PETD_01|08|SL|1|corr_file_size
0017|GEMS_PETD_01|09|LO|1|scan_id
0017|GEMS_PETD_01|0a|DT|1|scan_datetime
0017|GEMS_PETD_01|0b|LO|1|norm_2d_cal_id
0017|GEMS_PETD_01|0c|SH|1|hosp_identifier
0017|GEMS_PETD_01|0d|SL|1|archived
0019|GEMS_PETD_01|01|UI|1|wc_cal_id
0019|GEMS_PETD_01|02|SH|1|compatible_version
0019|GEMS_PETD_01|03|SH|1|software_version
0019|GEMS_PETD_01|04|DT|1|cal_datetime
0019|GEMS_PETD_01|05|SL|1|cal_type
0019|GEMS_PETD_01|06|LO|1|cal_description
0019|GEMS_PETD_01|07|LO|1|cal_hardware
0019|GEMS_PETD_01|08|OB|1|coefficients
0019|GEMS_PETD_01|0a|FL|1|activity_factor_hs
0019|GEMS_PETD_01|0b|FL|1|activity_factor_3d
0019|GEMS_PETD_01|0c|LO|1|scan_id
0019|GEMS_PETD_01|0d|DT|1|scan_datetime
0019|GEMS_PETD_01|0e|SH|1|hosp_identifier
0019|GEMS_PETD_01|0f|FL|1|meas_activity
0019|GEMS_PETD_01|10|DT|1|meas_datetime
0019|GEMS_PETD_01|11|SL|1|axial_filter_3d
0019|GEMS_PETD_01|12|FL|1|axial_cutoff_3d
0019|GEMS_PETD_01|13|SL|1|default_flag
0019|GEMS_PETD_01|14|SL|1|archived
0019|GEMS_PETD_01|15|SL|1|wc_cal_rec_method
0019|GEMS_PETD_01|16|SL|1|activity_factor_2d
0019|GEMS_PETD_01|17|SL|1|isotope
0021|GEMS_PETD_01|01|US|1|raw_data_type
0021|GEMS_PETD_01|02|UL|1|raw_data_size
5001|GEMS_PETD_01|02|SH|1|Curve Compatible Version
5001|GEMS_PETD_01|03|SH|1|Curve Software Version
5001|GEMS_PETD_01|04|SL|1|Statistics Type
5001|GEMS_PETD_01|05|LT|1|How Derived
5001|GEMS_PETD_01|06|SL|1|How Derived Size
5001|GEMS_PETD_01|07|SL|1|Multi Patient
5001|GEMS_PETD_01|08|SL|1|Deadtime
5003|GEMS_PETD_01|01|SQ|1|Graph Sequence
5003|GEMS_PETD_01|02|UI|1|Graph ID
5003|GEMS_PETD_01|03|SH|1|Graph Compatible Version
5003|GEMS_PETD_01|04|SH|1|Graph Software Version
5003|GEMS_PETD_01|05|LO|1|Title
5003|GEMS_PETD_01|06|DT|1|Graph Date Time
5003|GEMS_PETD_01|07|ST|1|Graph Description
5003|GEMS_PETD_01|08|LO|1|Title Font Name
5003|GEMS_PETD_01|09|SH|1|Title Font Size
5003|GEMS_PETD_01|0a|LO|1|Footer
5003|GEMS_PETD_01|0b|SH|1|Footer Font Size
5003|GEMS_PETD_01|0c|LO|1|Foreground Color
5003|GEMS_PETD_01|0d|LO|1|Background Color
5003|GEMS_PETD_01|0e|SL|1|Graph Border
5003|GEMS_PETD_01|0f|SL|1|Graph Width
5003|GEMS_PETD_01|10|SL|1|Graph Height
5003|GEMS_PETD_01|11|SL|1|Grid
5003|GEMS_PETD_01|12|LO|1|Label Font Name
5003|GEMS_PETD_01|13|SH|1|Label Font Size
5003|GEMS_PETD_01|14|LO|1|Axes Color
5003|GEMS_PETD_01|15|LO|1|X Axis Label
5003|GEMS_PETD_01|16|SL|1|X Axis Units
5003|GEMS_PETD_01|17|FL|1|X Major Tics
5003|GEMS_PETD_01|18|FL|1|X Axis Min
5003|GEMS_PETD_01|19|FL|1|X Axis Max
5003|GEMS_PETD_01|1a|LO|1|Y Axis Label
5003|GEMS_PETD_01|1b|SL|1|Y Axis Units
5003|GEMS_PETD_01|1c|FL|1|Y Major Tics
5003|GEMS_PETD_01|1d|FL|1|Y Axis Min
5003|GEMS_PETD_01|1e|FL|1|Y Axis Max
5003|GEMS_PETD_01|1f|LO|1|Legend Font Name
5003|GEMS_PETD_01|20|SH|1|Legend Font Size
5003|GEMS_PETD_01|21|SL|1|Legend Location X
5003|GEMS_PETD_01|22|SL|1|Legend Location Y
5003|GEMS_PETD_01|23|SL|1|Legend Width
5003|GEMS_PETD_01|24|SL|1|Legend Height
5003|GEMS_PETD_01|25|SL|1|Legend Border
5003|GEMS_PETD_01|26|SL|1|Multi Patient
5005|GEMS_PETD_01|01|SQ|1|Curve Presentation Sequence
5005|GEMS_PETD_01|02|UI|1|Curve Presentation ID
5005|GEMS_PETD_01|03|UI|1|Graph ID
5005|GEMS_PETD_01|04|UI|1|Curve ID
5005|GEMS_PETD_01|05|SH|1|Curve Presentation Compatible Version
5005|GEMS_PETD_01|06|SH|1|Curve Presentation Software Version
5005|GEMS_PETD_01|07|LO|1|Curve Label
5005|GEMS_PETD_01|08|LO|1|Color
5005|GEMS_PETD_01|09|SL|1|Line Type
5005|GEMS_PETD_01|0a|SL|1|Line Width
5005|GEMS_PETD_01|0b|SL|1|Point Symbol
5005|GEMS_PETD_01|0c|SL|1|Point Symbol Dim
5005|GEMS_PETD_01|0d|LO|1|Point Color
0009|GEMS_GENIE_1|01|SH|1|Unknown
0009|GEMS_GENIE_1|28|SL|1|Number RR Windows
0009|GEMS_GENIE_1|2b|LO|1|Trigger History UID
0009|GEMS_GENIE_1|2f|SL|1|Table Direction
0009|GEMS_GENIE_1|33|FD|1|Rotational Continuous Speed
0009|GEMS_GENIE_1|34|SL|1|Gantry Motion Type (Retired)
0009|GEMS_GENIE_1|44|SL|1|Num Views Acquired (Retired)
0009|GEMS_GENIE_1|45|LT|1|Unknown
0009|GEMS_GENIE_1|46|UI|1|Unknown
0011|GEMS_GENIE_1|11|SL|1|Dataset Modified
0011|GEMS_GENIE_1|14|LO|1|Completion Time
0011|GEMS_GENIE_1|1e|SL|4|Energy Width (Retired)
0011|GEMS_GENIE_1|21|DS|1|Acq Zoom (Retired)
0011|GEMS_GENIE_1|22|DS|1|Acq Pan (Retired)
0011|GEMS_GENIE_1|29|SL|1|Uniformity Mean
0011|GEMS_GENIE_1|2a|FD|1|Phase Duration (Retired)
0011|GEMS_GENIE_1|2c|FD|1|View X Adjustment
0011|GEMS_GENIE_1|2d|FD|1|View Y Adjustment
0011|GEMS_GENIE_1|2e|SL|1|Pixel Overflow Flag
0011|GEMS_GENIE_1|2f|SL|1|Overflow Level
0011|GEMS_GENIE_1|31|LO|1|Acquisition Parent UID
0011|GEMS_GENIE_1|32|LO|1|Processing Parent UID
0011|GEMS_GENIE_1|39|SL|1|Compression Type
0011|GEMS_GENIE_1|3d|SL|4|Energy Peak (Retired)
0011|GEMS_GENIE_1|40|LO|1|Viewing Object Name
0011|GEMS_GENIE_1|41|SL|1|Orientation Angle
0011|GEMS_GENIE_1|42|FD|1|Rotation Angle
0011|GEMS_GENIE_1|43|SL|1|Window Inverse Flag
0011|GEMS_GENIE_1|50|LO|1|Where Object Name
0011|GEMS_GENIE_1|57|FD|2|FOV
0011|GEMS_GENIE_1|61|SL|1|Image Size
0011|GEMS_GENIE_1|62|FD|1|Linear FOV
0011|GEMS_GENIE_1|63|FD|1|Spatial Offset
0011|GEMS_GENIE_1|64|FD|1|Spatial Orientation
0011|GEMS_GENIE_1|65|LO|1|Reference Dataset UID
0011|GEMS_GENIE_1|66|SH|1|Starcam Reference Dataset
0011|GEMS_GENIE_1|67|SL|1|Reference Frame Number
0011|GEMS_GENIE_1|68|SL|1|Cursor Length
0011|GEMS_GENIE_1|69|SL|1|Number of Cursors
0011|GEMS_GENIE_1|6a|SL|1|Cursor Coordinates
0011|GEMS_GENIE_1|6b|SL|1|Recon Options Flag
0011|GEMS_GENIE_1|6c|FD|1|Motion Threshold
0011|GEMS_GENIE_1|6d|UI|1|Motion Curve UID
0011|GEMS_GENIE_1|6e|SL|1|Recon Type
0011|GEMS_GENIE_1|6f|SL|1|Pre Filter Type
0011|GEMS_GENIE_1|71|SL|1|Back Proj Filter Type
0011|GEMS_GENIE_1|72|SL|1|Recon Arc
0011|GEMS_GENIE_1|73|FD|1|Recon Pan AP Offset
0011|GEMS_GENIE_1|74|FD|1|Recon Pan LR Offset
0011|GEMS_GENIE_1|75|FD|1|Recon Area
0011|GEMS_GENIE_1|76|SL|1|Start View
0011|GEMS_GENIE_1|77|SL|1|Attenuation Type
0011|GEMS_GENIE_1|78|SL|1|Dua lEnergy Processing
0011|GEMS_GENIE_1|79|SH|1|Pre Filter Param
0011|GEMS_GENIE_1|7a|SH|1|Pre Filter Param 2
0011|GEMS_GENIE_1|7b|SH|1|Back Proj Filter Param
0011|GEMS_GENIE_1|7c|SH|1|Back Proj Filter Param 2
0011|GEMS_GENIE_1|7d|SH|1|Attenuation Coef
0011|GEMS_GENIE_1|7e|SL|1|Ref Slice Width
0011|GEMS_GENIE_1|7f|FD|1|Ref Trans Pixel Volume
0011|GEMS_GENIE_1|81|SH|1|Attenuation Threshold
0011|GEMS_GENIE_1|82|FD|1|Interpolation Distance
0011|GEMS_GENIE_1|83|FD|1|Interpolation Center X
0011|GEMS_GENIE_1|84|FD|1|Interpolation Center Y
0011|GEMS_GENIE_1|85|SL|1|Quant Filter Flag
0011|GEMS_GENIE_1|86|SL|1|Head Conversion
0011|GEMS_GENIE_1|87|SL|1|Slice Width Pixels
0011|GEMS_GENIE_1|88|SL|1|Rfmtr Trans Ref
0011|GEMS_GENIE_1|89|FD|1|Rfmtr Trans Ref mm
0011|GEMS_GENIE_1|8a|SL|1|Two Line Trans Ref
0011|GEMS_GENIE_1|8b|SL|1|Three-D Zero
0011|GEMS_GENIE_1|8c|SL|1|Three-D Zero Length
0011|GEMS_GENIE_1|8d|SL|1|Three-D Zero In
0011|GEMS_DL_PATNT_01|80|UI|1|Patient Instance Uid
0011|GEMS_DL_PATNT_01|81|IS|1|Last Study Number
0011|GEMS_DL_PATNT_01|82|CS|1|Patient Repaired
0011|GEMS_DL_PATNT_01|83|CS|1|Lock Demographics
0013|GEMS_GENIE_1|13|SQ|1|eNTEGRA Frame Sequence
0013|GEMS_GENIE_1|14|SL|1|Original Image Number
0013|GEMS_GENIE_1|15|FD|1|Fscalar
0013|GEMS_GENIE_1|1b|FD|1|Det Ang Separation
0013|GEMS_GENIE_1|20|FD|1|Accepted Beats Time
0013|GEMS_GENIE_1|21|FD|2|Threshold
0013|GEMS_GENIE_1|22|FD|2|Linear Depth
0013|GEMS_GENIE_1|23|LO|1|Unif Date Time
0013|GEMS_GENIE_1|24|SL|1|Series Accepted Beats
0013|GEMS_GENIE_1|25|SL|1|Series Rejected Beats
0015|GEMS_GENIE_1|10|SL|1|Frame Termination Condition
0015|GEMS_GENIE_1|11|SL|1|Frame Termination Value
0015|GEMS_GENIE_1|12|SL|1|Num ECT Phases
0015|GEMS_GENIE_1|13|SL|1|Num WB Scans
0015|GEMS_GENIE_1|14|SL|1|ECT Phase Num
0015|GEMS_GENIE_1|15|SL|1|WB Scan Num
0015|GEMS_GENIE_1|16|SL|1|Comb Head Number
0015|GEMS_GENIE_1|17|UL|1|Preceding Beat
0015|GEMS_DL_STUDY_01|80|DS|1|Study Dose
0015|GEMS_DL_STUDY_01|81|DS|1|Study Total Dap
0015|GEMS_DL_STUDY_01|82|DS|1|Fluoro Dose Area Product
0015|GEMS_DL_STUDY_01|83|IS|1|Study Fluoro Time
0015|GEMS_DL_STUDY_01|84|DS|1|Cine Dose Area Product
0015|GEMS_DL_STUDY_01|85|IS|1|Study Record Time
0015|GEMS_DL_STUDY_01|86|IS|1|Last XA Number
0015|GEMS_DL_STUDY_01|88|PN|1-n|Def Operator Name
0015|GEMS_DL_STUDY_01|89|PN|1-n|Def Performing Physician Name
0015|GEMS_DL_STUDY_01|8a|CS|2|Def Patient Orientation
0015|GEMS_DL_STUDY_01|8b|IS|1|Last Sc Number
0015|GEMS_DL_STUDY_01|8e|UI|1|Common Series Instance UID
0015|GEMS_DL_STUDY_01|8f|IS|1|Study Number
0015|GEMS_DL_STUDY_01|92|FL|1|Unknown
0015|GEMS_DL_STUDY_01|93|FL|1|Unknown
0015|GEMS_DL_STUDY_01|94|FL|1|Unknown
0015|GEMS_DL_STUDY_01|95|IS|1|Unknown
0015|GEMS_DL_STUDY_01|96|FL|1|Unknown
0015|GEMS_DL_STUDY_01|97|IS|1|Unknown
0015|GEMS_DL_STUDY_01|98|FL|1|Unknown
0015|GEMS_DL_STUDY_01|99|FL|1|Unknown
0015|GEMS_DL_STUDY_01|9a|FL|1|Unknown
0015|GEMS_DL_STUDY_01|9b|IS|1|Unknown
0015|GEMS_DL_STUDY_01|9c|FL|1|Unknown
0015|GEMS_DL_STUDY_01|9d|IS|1|Unknown
0015|GEMS_DL_SERIES_01|85|LO|1|Series File Name
0015|GEMS_DL_SERIES_01|87|IS|1|Number of Images
0015|GEMS_DL_SERIES_01|8c|CS|1|Sent Flag
0015|GEMS_DL_SERIES_01|8d|US|1|Item Locked
0019|GEMS_GENIE_1|5f|SQ|1|Unknown
0019|GEMS_DL_IMG_01|0b|DS|40909|FOV Dimension Double
0019|GEMS_DL_IMG_01|2b|FL|1|Distance to table top
0019|GEMS_DL_IMG_01|30|LO|1|Image File Name
0019|GEMS_DL_IMG_01|31|IS|1|Default Spatial Filter Family
0019|GEMS_DL_IMG_01|32|IS|1|Default Spatial Filter Strength
0019|GEMS_DL_IMG_01|33|DS|1|Min Saturation Dose
0019|GEMS_DL_IMG_01|34|DS|1|Detector Gain
0019|GEMS_DL_IMG_01|35|DS|1|Patient Dose Limit
0019|GEMS_DL_IMG_01|36|DS|1|Preproc Image Rate Max
0019|GEMS_DL_IMG_01|37|CS|1|Sensor Roi Shape
0019|GEMS_DL_IMG_01|38|DS|1|Sensor Roi x Position
0019|GEMS_DL_IMG_01|39|DS|1|Sensor Roi y Position
0019|GEMS_DL_IMG_01|3a|DS|1|Sensor Roi x Size
0019|GEMS_DL_IMG_01|3b|DS|1|Sensor Roi y Size
0019|GEMS_DL_IMG_01|3d|DS|1|Noise Sensitivity
0019|GEMS_DL_IMG_01|3e|DS|1|Sharp Sensitivity
0019|GEMS_DL_IMG_01|3f|DS|1|Contrast Sensitivity
0019|GEMS_DL_IMG_01|40|DS|1|Lag Sensitivity
0019|GEMS_DL_IMG_01|41|CS|1|Tube
0019|GEMS_DL_IMG_01|42|US|1|Detector Size Rows
0019|GEMS_DL_IMG_01|43|US|1|Detector Size Columns
0019|GEMS_DL_IMG_01|44|DS|1|Min Object Size
0019|GEMS_DL_IMG_01|45|DS|1|Max Object Size
0019|GEMS_DL_IMG_01|46|DS|1|Max Object Speed
0019|GEMS_DL_IMG_01|47|CS|1|Object Back Motion
0019|GEMS_DL_IMG_01|48|UL|1|Exposure Trajectory Family
0019|GEMS_DL_IMG_01|49|DS|1|Window Time Duration
0019|GEMS_DL_IMG_01|4a|CS|1|Positioner Angle Display Mode
0019|GEMS_DL_IMG_01|4b|IS|2|Detector Origin
0019|GEMS_DL_IMG_01|4c|CS|1|Unknown
0019|GEMS_DL_IMG_01|4e|DS|2|Default Brightness and Contrast
0019|GEMS_DL_IMG_01|4f|DS|2|User Brightness and Contrast
0019|GEMS_DL_IMG_01|50|IS|1|Source Series Number
0019|GEMS_DL_IMG_01|51|IS|1|Source Image Number
0019|GEMS_DL_IMG_01|52|IS|1|Source Frame Number
0019|GEMS_DL_IMG_01|53|UI|1|Source Series Item Id
0019|GEMS_DL_IMG_01|54|UI|1|Source Image Item Id
0019|GEMS_DL_IMG_01|55|UI|1|Source Frame Item Id
0019|GEMS_DL_IMG_01|60|US|1|Number of Points Before Acquisition
0019|GEMS_DL_IMG_01|61|OW|1|Curve Data Before Acquisition
0019|GEMS_DL_IMG_01|62|US|1|Number of Points Trigger
0019|GEMS_DL_IMG_01|63|OW|1|Curve Data Trigger
0019|GEMS_DL_IMG_01|64|SH|1|ECG Synchronization
0019|GEMS_DL_IMG_01|65|SH|1|ECG Delay Mode
0019|GEMS_DL_IMG_01|66|IS|1-n|ECG Delay Vector
0019|GEMS_DL_IMG_01|67|DS|1|Unknown
0019|GEMS_DL_IMG_01|68|DS|1|Unknown
0019|GEMS_DL_IMG_01|69|DS|1|Unknown
0019|GEMS_DL_IMG_01|7a|DS|1|Unknown
0019|GEMS_DL_IMG_01|7b|DS|1|Unknown
0019|GEMS_DL_IMG_01|7c|DS|1|Unknown
0019|GEMS_DL_IMG_01|80|DS|1|Image Dose
0019|GEMS_DL_IMG_01|81|US|1|Calibration Frame
0019|GEMS_DL_IMG_01|82|CS|1|Calibration Object
0019|GEMS_DL_IMG_01|83|DS|1|Calibration Object Size mm
0019|GEMS_DL_IMG_01|84|FL|1|Calibration Factor
0019|GEMS_DL_IMG_01|85|DA|1|Calibration Date
0019|GEMS_DL_IMG_01|86|TM|1|Calibration Time
0019|GEMS_DL_IMG_01|87|US|1|Calibration Accuracy
0019|GEMS_DL_IMG_01|88|CS|1|Calibration Extended
0019|GEMS_DL_IMG_01|89|US|1|Calibration Image Original
0019|GEMS_DL_IMG_01|8a|US|1|Calibration Frame Original
0019|GEMS_DL_IMG_01|8b|US|1|Calibration nb points uif
0019|GEMS_DL_IMG_01|8c|US|1-n|Calibration Points Row
0019|GEMS_DL_IMG_01|8d|US|1-n|Calibration Points Column
0019|GEMS_DL_IMG_01|8e|FL|1|Calibration Magnification Ratio
0019|GEMS_DL_IMG_01|8f|LO|1|Calibration Software Version
0019|GEMS_DL_IMG_01|90|LO|1|Extended Calibration Software Version
0019|GEMS_DL_IMG_01|91|IS|1|Calibration Return Code
0019|GEMS_DL_IMG_01|92|DS|1|Detector Rotation Angle
0019|GEMS_DL_IMG_01|93|CS|1|Spatial Change
0019|GEMS_DL_IMG_01|94|CS|1|Inconsistent Flag
0019|GEMS_DL_IMG_01|95|CS|2|Horizontal and Vertical Image Flip
0019|GEMS_DL_IMG_01|96|CS|1|Internal Label Image
0019|GEMS_DL_IMG_01|97|DS|1-n|Angle 1 increment
0019|GEMS_DL_IMG_01|98|DS|1-n|Angle 2 increment
0019|GEMS_DL_IMG_01|99|DS|1-n|Angle 3 increment
0019|GEMS_DL_IMG_01|9a|DS|1-n|Sensor Feedback
0019|GEMS_DL_IMG_01|9b|CS|1|Grid
0019|GEMS_DL_IMG_01|9c|FL|1|Default Mask Pixel Shift
0019|GEMS_DL_IMG_01|9d|CS|1|Applicable Review Mode
0019|GEMS_DL_IMG_01|9e|DS|1-n|Log LUT Control Points
0019|GEMS_DL_IMG_01|9f|DS|1-n|Exp LUT SUB Control Points
0019|GEMS_DL_IMG_01|a0|DS|1|ABD Value
0019|GEMS_DL_IMG_01|a1|DS|1|Subtraction Window Center
0019|GEMS_DL_IMG_01|a2|DS|1|Subtraction Window Width
0019|GEMS_DL_IMG_01|a3|DS|1|Image Rotation
0019|GEMS_DL_IMG_01|a4|CS|1|Auto Injection Enabled
0019|GEMS_DL_IMG_01|a5|CS|1|Injection Phase
0019|GEMS_DL_IMG_01|a6|DS|1|Injection Delay
0019|GEMS_DL_IMG_01|a7|IS|1|Reference Injection Frame Number
0019|GEMS_DL_IMG_01|a8|DS|1|Injection Duration
0019|GEMS_DL_IMG_01|a9|DS|1-n|EPT
0019|GEMS_DL_IMG_01|aa|CS|1|Can Downscan 512
0019|GEMS_DL_IMG_01|ab|IS|1|Current Spatial Filter Strength
0019|GEMS_DL_IMG_01|ac|DS|1|Brightness Sensitivity
0019|GEMS_DL_IMG_01|ad|DS|1-n|Exp LUT NOSUB Control Points
0019|GEMS_DL_IMG_01|af|DS|1-n|Unknown
0019|GEMS_DL_IMG_01|b0|DS|1-n|Unknown
0019|GEMS_DL_IMG_01|b1|LO|1|Acquisition Mode Description
0019|GEMS_DL_IMG_01|b2|LO|1|Acquisition Mode Description Label
0019|GEMS_DL_IMG_01|b3|LO|1|Unknown
0019|GEMS_DL_IMG_01|b8|FL|1|Unknown
0019|GEMS_DL_IMG_01|ba|CS|1|Acquisition Region
0019|GEMS_DL_IMG_01|bb|CS|1|Acquisition SUB Mode
0019|GEMS_DL_IMG_01|bc|FL|1|Table Cradle Angle
0019|GEMS_DL_IMG_01|bd|CS|1-n|Table Rotation Status Vector
0019|GEMS_DL_IMG_01|be|FL|1-n|Source to Image Distance per Frame Vector
0019|GEMS_DL_IMG_01|c2|DS|1-n|Unknown
0019|GEMS_DL_IMG_01|c3|FL|1-n|Table Rotation Angle Increment
0019|GEMS_DL_IMG_01|c4|IS|1|Unknown
0019|GEMS_DL_IMG_01|c7|CS|1|Patient Position per Image
0019|GEMS_DL_IMG_01|d7|FL|1-n|Table X Position to Iso‐center Increment
0019|GEMS_DL_IMG_01|d8|FL|1-n|Table Y Position to Iso‐center Increment
0019|GEMS_DL_IMG_01|d9|FL|1-n|Table Z Position to Iso‐center Increment
0019|GEMS_DL_IMG_01|da|FL|1-n|Table Head Tilt Angle Increment
0019|GEMS_DL_IMG_01|dc|LO|1|Unknown
0019|GEMS_DL_IMG_01|de|CS|1|Acquisition Plane
0019|GEMS_DL_IMG_01|dd|DS|1|Unknown
0019|GEMS_DL_IMG_01|e0|FL|1|Unknown
0019|GEMS_DL_IMG_01|e9|FL|1-n|Source to Detector Distance per Frame Vector
0019|GEMS_DL_IMG_01|ea|FL|1|Table Rotation Angle
0019|GEMS_DL_IMG_01|eb|FL|1|Table X Position to Iso‐center
0019|GEMS_DL_IMG_01|ec|FL|1|Table Y Position to Iso‐center
0019|GEMS_DL_IMG_01|ed|FL|1|Table Z Position to Iso‐center
0019|GEMS_DL_IMG_01|ee|FL|1|Table Head Tilt Angle
0019|GEMS_DL_IMG_01|ef|FL|1|Unknown
0019|DLX_SERIE_01|20|LO|1|Ip Address
0019|DLX_SERIE_01|21|DS|1|Table position Z (vertical) first frame
0019|DLX_SERIE_01|22|DS|1|Table position X (longitudinal) first frame
0019|DLX_SERIE_01|23|DS|1|Table position Y (lateral) first frame
0019|DLX_SERIE_01|24|DS|1|Lambda cm Pincushion Distortion
0019|DLX_SERIE_01|25|DS|1|LV Regression Slope Coefficient
0019|DLX_SERIE_01|26|DS|1|LV Regression Intercept Coefficient
0019|DLX_SERIE_01|27|DS|1|Image chain FWHM psf mm min
0019|DLX_SERIE_01|28|DS|1|Image chain FWHM psf mm max
0019|GEMS_DL_SERIES_01|4c|CS|1|Internal Label
0019|GEMS_DL_SERIES_01|4d|CS|1|Browser Hide
0021|GEMS_XR3DCAL_01|20|LT|1|Generalized Calibration
0021|Mayo/IBM Archive Project|01|UN|1|Unknown
0021|Mayo/IBM Archive Project|10|UN|1|Unknown
0021|Mayo/IBM Archive Project|11|UN|1|Unknown
0021|Mayo/IBM Archive Project|12|UN|1|Unknown
0021|Mayo/IBM Archive Project|13|UN|1|Unknown
0021|Mayo/IBM Archive Project|14|UN|1|Unknown
0021|Mayo/IBM Archive Project|15|UN|1|Unknown
0021|Mayo/IBM Archive Project|16|UN|1|Unknown
0021|Mayo/IBM Archive Project|17|UN|1|Unknown
0021|Mayo/IBM Archive Project|18|UN|1|Unknown
0021|Mayo/IBM Archive Project|19|UN|1|Unknown
0021|Mayo/IBM Archive Project|1a|UN|1|Unknown
0021|Mayo/IBM Archive Project|1b|UN|1|Unknown
0021|Mayo/IBM Archive Project|1c|UN|1|Unknown
0021|Mayo/IBM Archive Project|1d|UN|1|Unknown
0021|Mayo/IBM Archive Project|1e|UN|1|Unknown
0021|Mayo/IBM Archive Project|1f|UN|1|Unknown
0021|Mayo/IBM Archive Project|20|UN|1|Unknown
0021|Mayo/IBM Archive Project|40|UN|1|Unknown
0021|Mayo/IBM Archive Project|41|UN|1|Unknown
0021|Mayo/IBM Archive Project|50|UN|1|Unknown
0021|Mayo/IBM Archive Project|60|UN|1|Unknown
0021|Mayo/IBM Archive Project|65|UN|1|Unknown
0023|GEMS_3D_INTVL_01|01|SQ|1|X-Ray Marker Sequence
0023|GEMS_3D_INTVL_01|02|SH|1|Marker ID
0023|GEMS_3D_INTVL_01|03|CS|1|Marker Type
0023|GEMS_3D_INTVL_01|04|FL|1|Marker Size
0023|GEMS_3D_INTVL_01|05|US|3|Marker Color CIELab Value
0023|GEMS_3D_INTVL_01|06|LO|1|Marker Label
0023|GEMS_3D_INTVL_01|07|CS|1|Marker Visible State
0023|GEMS_3D_INTVL_01|08|LO|1|Marker Description
0023|GEMS_3D_INTVL_01|10|SQ|1|Marker Points Sequence
0023|GEMS_3D_INTVL_01|11|SH|1|Marker Point ID
0023|GEMS_3D_INTVL_01|12|FL|3|Marker Point Position
0023|GEMS_3D_INTVL_01|13|FL|1|Marker Point Size
0023|GEMS_3D_INTVL_01|14|US|3|Marker Point Color CIELab Value
0023|GEMS_3D_INTVL_01|16|CS|1|Marker Point Visible State
0023|GEMS_3D_INTVL_01|17|IS|1|Marker Point Order
0023|GEMS_3D_INTVL_01|18|FL|3|Volume Manual Registration
0023|GEMS_3D_INTVL_01|20|IS|1-n|Volumes Threshold
0023|GEMS_3D_INTVL_01|25|CS|1|Cut Plane Activation Flag
0023|GEMS_3D_INTVL_01|26|IS|1|Cut Plane Position Value
0023|GEMS_3D_INTVL_01|27|FL|3|Cut Plane Normal Value
0023|GEMS_3D_INTVL_01|28|FL|1|Volume Scaling Factor
0023|GEMS_3D_INTVL_01|29|FL|1|ROI to Table Top Distance
0023|GEMS_3D_INTVL_01|30|IS|1-n|DRR Threshold
0023|GEMS_3D_INTVL_01|31|FL|3|Volume Table Position
0023|GEMS_3D_INTVL_01|32|IS|1|Rendering Mode
0023|GEMS_3D_INTVL_01|33|IS|1|3D Object Opacity
0023|GEMS_3D_INTVL_01|34|IS|1|Invert Image
0023|GEMS_3D_INTVL_01|35|IS|1|Enhance Full
0023|GEMS_3D_INTVL_01|36|FL|1|Zoom
0023|GEMS_3D_INTVL_01|37|IS|2|Roam
0023|GEMS_3D_INTVL_01|38|IS|1|Window Level
0023|GEMS_3D_INTVL_01|39|IS|1|Window Width
0023|GEMS_3D_INTVL_01|40|CS|1|BMC Setting
0023|GEMS_3D_INTVL_01|41|CS|1|Back View Setting
0023|GEMS_3D_INTVL_01|42|CS|1-n|Sub Volume Visibility
0023|GEMS_3D_INTVL_01|43|CS|1|3D Landmarks Visibility
0023|GEMS_3D_INTVL_01|44|CS|1|Ablation Point Visibility
0025|GEMS_DL_FRAME_01|02|IS|1|Frame ID
0025|GEMS_DL_FRAME_01|03|DS|1|Distance Source to Detector
0025|GEMS_DL_FRAME_01|04|DS|1|Distance Source to Patient
0025|GEMS_DL_FRAME_01|05|DS|1|Distance Source to Skin
0025|GEMS_DL_FRAME_01|06|DS|1|Positioner Primary Angle
0025|GEMS_DL_FRAME_01|07|DS|1|Positioner Secondary Angle
0025|GEMS_DL_FRAME_01|08|IS|1|Beam Orientation
0025|GEMS_DL_FRAME_01|09|DS|1|L Arm Angle
0025|GEMS_DL_FRAME_01|0a|SQ|1|Frame Sequence
0025|GEMS_SERS_01|1b|OB|1|Protocol Data Block (compressed)
0025|GEMS_DL_FRAME_01|10|DS|1|Pivot Angle
0025|GEMS_DL_FRAME_01|1a|DS|1|Arc Angle
0025|GEMS_DL_FRAME_01|1b|DS|1|Table Vertical Position
0025|GEMS_DL_FRAME_01|1c|DS|1|Table Longitudinal Position
0025|GEMS_DL_FRAME_01|1d|DS|1|Table Lateral Position
0025|GEMS_DL_FRAME_01|1e|IS|1|Beam Cover Area
0025|GEMS_DL_FRAME_01|1f|DS|1|kVP Actual
0025|GEMS_DL_FRAME_01|20|DS|1|mAS Actual
0025|GEMS_DL_FRAME_01|21|DS|1|PW Actual
0025|GEMS_DL_FRAME_01|22|DS|1|Kvp Commanded
0025|GEMS_DL_FRAME_01|23|DS|1|Mas Commanded
0025|GEMS_DL_FRAME_01|24|DS|1|Pw Commanded
0025|GEMS_DL_FRAME_01|25|CS|1|Grid
0025|GEMS_DL_FRAME_01|26|DS|1|Sensor Feedback
0025|GEMS_DL_FRAME_01|27|DS|1|Target Entrance Dose
0025|GEMS_DL_FRAME_01|28|DS|1|Cnr Commanded
0025|GEMS_DL_FRAME_01|29|DS|1|Contrast Commanded
0025|GEMS_DL_FRAME_01|2a|DS|1|EPT Actual
0025|GEMS_DL_FRAME_01|2b|IS|1|Spectral Filter Znb
0025|GEMS_DL_FRAME_01|2c|DS|1|Spectral Filter Weight
0025|GEMS_DL_FRAME_01|2d|DS|1|Spectral Filter Density
0025|GEMS_DL_FRAME_01|2e|IS|1|Spectral Filter Thickness
0025|GEMS_DL_FRAME_01|2f|IS|1|Spectral Filter Status
0025|GEMS_DL_FRAME_01|30|IS|2|FOV Dimension
0025|GEMS_DL_FRAME_01|33|IS|2|FOV Origin
0025|GEMS_DL_FRAME_01|34|IS|1|Collimator Left Vertical Edge
0025|GEMS_DL_FRAME_01|35|IS|1|Collimator Right Vertical Edge
0025|GEMS_DL_FRAME_01|36|IS|1|Collimator Up Horizontal Edge
0025|GEMS_DL_FRAME_01|37|IS|1|Collimator Low Horizontal Edge
0025|GEMS_DL_FRAME_01|38|IS|1|Vertices Polygonal Collimator
0025|GEMS_DL_FRAME_01|39|IS|1|Contour Filter Distance
0025|GEMS_DL_FRAME_01|3a|UL|1|Contour Filter Angle
0025|GEMS_DL_FRAME_01|3b|CS|1|Table Rotation Status
0025|GEMS_DL_FRAME_01|3c|CS|1|Internal Label Frame
0033|GEMS_GENIE_1|07|LO|1-n|Original SOP Instance UID
0033|GEMS_GENIE_1|08|CS|1|eNTEGRA Data Object Type
0033|GEMS_GENIE_1|10|SL|1|Modified
0033|GEMS_GENIE_1|11|LO|1|Name
0033|GEMS_GENIE_1|16|LO|1|Protocol Data UID
0033|GEMS_GENIE_1|17|SH|1|Date
0033|GEMS_GENIE_1|18|SH|1|Time
0033|GEMS_GENIE_1|19|UL|1|Protocol Data Flags
0033|GEMS_GENIE_1|1a|UL|1|Protocol Name
0033|GEMS_GENIE_1|1b|LO|1|Relevant Data UID
0033|GEMS_GENIE_1|1c|LO|1|Bulk Data
0033|GEMS_GENIE_1|1d|SL|1-n|Int Data
0033|GEMS_GENIE_1|1e|FD|1-n|Double Data
0033|GEMS_GENIE_1|1f|OB|1|String Data
0033|GEMS_GENIE_1|20|LT|1-n|Bulk Data Format
0033|GEMS_GENIE_1|21|LT|1-n|Int Data Format
0033|GEMS_GENIE_1|22|LT|1-n|Double Data Format
0033|GEMS_GENIE_1|23|LT|1-n|String Data Format
0033|GEMS_GENIE_1|24|LT|1|Description
0033|GEMS_GENIE_1|30|UL|1|Allocate Trigger Buffer
0033|GEMS_GENIE_1|33|UL|1|Number of Triggers
0033|GEMS_GENIE_1|34|UL|1|Trigger Size
0033|GEMS_GENIE_1|35|UL|1|Trigger Data Size
0033|GEMS_GENIE_1|36|OB|1|Trigger Data
0035|GEMS_GENIE_1|01|FD|1-n|Start Angle
0039|GEMS_ADWSoft_DPO|aa|CS|1|Private Entity Type
0039|GEMS_ADWSoft_DPO1|95|LO|1|Unknown
0039|GEMS_AWSoft_SB1|50|UI|1|Reference to Study UID
0039|GEMS_AWSoft_SB1|51|UI|1|Reference to Series UID
0039|GEMS_AWSoft_SB1|52|IS|1|Reference to Original Instance Number
0039|GEMS_AWSoft_SB1|95|LO|1|Private Entity Launch Command
0039|GEMS_AWSOFT_CD1|65|UI|1|Reference to Study UID
0039|GEMS_AWSOFT_CD1|70|UI|1|Reference to Series UID
0039|GEMS_AWSOFT_CD1|75|IS|1|Reference to Original Instance Number
0039|GEMS_AWSOFT_CD1|80|IS|1|DPO Number
0039|GEMS_AWSOFT_CD1|85|DA|1|DPO Date
0039|GEMS_AWSOFT_CD1|90|TM|1|DPO Time
0039|GEMS_AWSOFT_CD1|95|LO|1|DPO Invocation String
0039|GEMS_AWSOFT_CD1|aa|CS|1|DPO Type
0039|GEMS_AWSOFT_CD1|ff|OB|1|DPO Data
0119|MRSC|11a5|DS|1-n|PhantRefValues
0043|GEMS_PARM_01|64|CS|1-n|Image Filter
0043|GEMS_PARM_01|66|US|1|Helical Correction Indicator
0043|GEMS_PARM_01|67|US|1|IBO Correction Indicator
0043|GEMS_PARM_01|68|US|1|XT Correction Indicator
0043|GEMS_PARM_01|69|US|1|Q-cal Correction Indicator
0043|GEMS_PARM_01|6a|US|1|AV Correction Indicator
0043|GEMS_PARM_01|6b|US|1|L-MDK Correction Indicator
0043|GEMS_PARM_01|6c|IS|1|Detector Row
0043|GEMS_PARM_01|6d|US|1|Area Size
0043|GEMS_PARM_01|6e|SH|1|Auto mA Mode
0043|GEMS_PARM_01|70|LO|1|Paradigm Name
0043|GEMS_PARM_01|71|ST|1|Paradigm Description
0043|GEMS_PARM_01|72|UI|1|Paradigm UID
0043|GEMS_PARM_01|73|US|1|Experiment Type
0043|GEMS_PARM_01|74|US|1|Number of Rest Volumes
0043|GEMS_PARM_01|75|US|1|Number of Active Volumes
0043|GEMS_PARM_01|76|US|1|Number of Dummy Scans
0043|GEMS_PARM_01|77|SH|1|Application Name
0043|GEMS_PARM_01|78|SH|1|Application Version
0043|GEMS_PARM_01|79|US|1|Slices Per Volume
0043|GEMS_PARM_01|7a|US|1|Expected Time Points
0043|GEMS_PARM_01|7b|FL|1-n|Regressor Values
0043|GEMS_PARM_01|7c|FL|1|Delay After Slice Group
0043|GEMS_PARM_01|7d|US|1|Recon Mode Flag Word
0043|GEMS_PARM_01|7e|LO|1-n|PACC Specific Information
0043|GEMS_PARM_01|7f|DS|1-n|Reserved
0043|GEMS_PARM_01|80|LO|1-n|Coil ID Data
0043|GEMS_PARM_01|81|LO|1|GE Coil Name
0043|GEMS_PARM_01|83|DS|40909|Asset R Factors
0043|GEMS_PARM_01|84|LO|5|Additional Asset Data
0043|GEMS_PARM_01|85|UT|1|Debug Data (Text Format)
0043|GEMS_PARM_01|86|OB|1|Debug Data (Binary Format)
0043|GEMS_PARM_01|87|UT|1|Reserved
0043|GEMS_PARM_01|88|UI|1|PURE Acquisition Calibration Series UID
0043|GEMS_PARM_01|89|LO|3|Governing Body, dB/dt, and SAR definition
0043|GEMS_PARM_01|8a|CS|1|Private In-Plane Phase Encoding Direction
0119|MRSC|1200|IS|1-n|ImageProcessStatus
0045|GEMS_SENO_02|1b|LO|1|Clinical View
0045|GEMS_SENO_02|1d|DS|1|Mean Of Raw Gray Levels
0045|GEMS_SENO_02|1e|DS|1|Mean Of Offset Gray Levels
0045|GEMS_SENO_02|1f|DS|1|Mean Of Corrected Gray Levels
0045|GEMS_SENO_02|49|DS|1|Radiological Thickness
0045|GEMS_SENO_02|50|UI|1|Fallback Instance UID (CR or SC)
0045|GEMS_SENO_02|51|UI|1|Fallback Series UID (CR or SC)
0045|GEMS_SENO_02|52|IS|1|Raw Diagnostic Low
0045|GEMS_SENO_02|53|IS|1|Raw Diagnostic High
0045|GEMS_SENO_02|54|DS|1|Exponent
0045|GEMS_SENO_02|55|IS|1|A Coefficients
0045|GEMS_SENO_02|56|DS|1|Noise Reduction Sensitivity
0045|GEMS_SENO_02|57|DS|1|Noise Reduction Threshold
0045|GEMS_SENO_02|58|DS|1|Mu
0045|GEMS_SENO_02|59|IS|1|Threshold
0045|GEMS_SENO_02|60|IS|4|Breast ROI X
0045|GEMS_SENO_02|61|IS|4|Breast ROI Y
0045|GEMS_SENO_02|62|IS|1|User Window Center
0045|GEMS_SENO_02|63|IS|1|User Window Width
0045|GEMS_SENO_02|64|IS|1|Segmentation Threshold
0045|GEMS_SENO_02|65|IS|1|Detector Entrance Dose
0045|GEMS_SENO_02|66|IS|1|Asymmetrical Collimation Information
0045|GEMS_SENO_02|71|OB|1|STX Buffer
0045|GEMS_SENO_02|72|DS|2|Image Crop Point
0045|GEMS_SENO_02|90|SH|1|Premium View Beta
0045|GEMS_SENO_02|a0|DS|1|Signal Average Factor
0045|GEMS_SENO_02|a1|DS|2-n|Organ Dose for Source Images
0045|GEMS_SENO_02|a2|DS|2-n|Entrance dose in mGy for Source Images
0045|GEMS_SENO_02|a4|DS|1|Organ Dose in dGy for Complete DBT Sequence
0045|GEMS_SENO_02|a6|UI|1|SOP Instance UID for Lossy Compression
0045|GEMS_SENO_02|a7|LT|1|Reconstruction Parameters
0045|GEMS_SENO_02|a8|DS|1|Entrance Dose in dGy for Complete DBT Sequence
0043|GEMS_PARM_01|8c|DS|1|Voxel Location
0043|GEMS_PARM_01|8d|DS|1-n|SAT Band Locations
0043|GEMS_PARM_01|8e|DS|3|Spectro Prescan Values
0043|GEMS_PARM_01|8f|DS|3|Spectro Parameters
0043|GEMS_PARM_01|90|LO|1-n|SAR Definition
0043|GEMS_PARM_01|91|DS|1-n|SAR Value
0043|GEMS_PARM_01|92|LO|1|Image Error Text
0043|GEMS_PARM_01|93|DS|1-n|Spectro Quantitation Values
0043|GEMS_PARM_01|94|DS|1-n|Spectro Ratio Values
0043|GEMS_PARM_01|95|LO|1|Prescan Reuse String
0043|GEMS_PARM_01|96|CS|1|Content Qualification
0043|GEMS_PARM_01|98|UI|1|ASSET Acquisition Calibration Series UID
0043|GEMS_PARM_01|99|LO|1-n|Extended Options
0043|GEMS_PARM_01|9a|IS|1|Rx Stack Identification
0045|GEMS_HELIOS_01|01|SS|1|Number of Macro Rows in Detector
0045|GEMS_HELIOS_01|02|FL|1|Macro width at ISO Center
0045|GEMS_HELIOS_01|03|SS|1|DAS type
0045|GEMS_HELIOS_01|04|SS|1|DAS gain
0045|GEMS_HELIOS_01|05|SS|1|DAS Temprature
0045|GEMS_HELIOS_01|06|CS|1|Table Direction
0045|GEMS_HELIOS_01|07|FL|1|Z smoothing Factor
0045|GEMS_HELIOS_01|08|SS|1|View Weighting Mode
0045|GEMS_HELIOS_01|09|SS|1|Sigma Row number
0047|GEMS_ADWSoft_3D1|8a|US|1|Number Of Injections
0047|GEMS_ADWSoft_3D1|8b|US|1|Frame Count
0047|GEMS_ADWSoft_3D1|9a|DS|9|Transform Rotation Matrix
0047|GEMS_ADWSoft_3D1|9b|DS|3|Transform Translation Vector
0047|GEMS_ADWSoft_3D1|9c|LO|1|Transform Label
0047|GEMS_ADWSoft_3D1|b0|SQ|1|Wireframe List
0047|GEMS_ADWSoft_3D1|b1|US|1|Wireframe Count
0047|GEMS_ADWSoft_3D1|b2|US|1|Location System
0047|GEMS_ADWSoft_3D1|b5|LO|1|Wireframe Name
0047|GEMS_ADWSoft_3D1|b6|LO|1|Wireframe Group Name
0047|GEMS_ADWSoft_3D1|b7|LO|1|Wireframe Color
0047|GEMS_ADWSoft_3D1|b8|SL|1|Wireframe Attributes
0047|GEMS_ADWSoft_3D1|b9|SL|1|Wireframe Point Count
0047|GEMS_ADWSoft_3D1|ba|SL|1|Wireframe Timestamp
0047|GEMS_ADWSoft_3D1|bb|SQ|1|Wireframe Point List
0047|GEMS_ADWSoft_3D1|bc|DS|3|Wireframe Points Coordinates
0047|GEMS_ADWSoft_3D1|c0|DS|3|Volume Upper Left High Corner RAS
0047|GEMS_ADWSoft_3D1|c1|DS|9|Volume Slice To RAS Rotation Matrix
0047|GEMS_ADWSoft_3D1|c2|DS|1|Volume Upper Left High Corner TLOC
0047|GEMS_ADWSoft_3D1|d1|OB|1|Volume Segment List
0047|GEMS_ADWSoft_3D1|d2|OB|1|Volume Gradient List
0047|GEMS_ADWSoft_3D1|d3|OB|1|Volume Density List
0047|GEMS_ADWSoft_3D1|d4|OB|1|Volume Z Position List
0047|GEMS_ADWSoft_3D1|d5|OB|1|Volume Original Index List
0047|GEMS_3DSTATE_001|e9|FL|3|Unknown
0047|GEMS_3DSTATE_001|ea|DS|3|Unknown
0047|GEMS_3DSTATE_001|eb|DS|3|Unknown
0047|GEMS_3DSTATE_001|ec|FL|1|Unknown
0047|GEMS_3DSTATE_001|ed|CS|1|Unknown
0045|GEMS_HELIOS_01|0b|FL|1|Maximum Offset Value
0045|GEMS_HELIOS_01|0c|SS|1|Number of Views shifted
0045|GEMS_HELIOS_01|0d|SS|1|Z tracking Flag
0045|GEMS_HELIOS_01|0e|FL|1|Mean Z error
0045|GEMS_HELIOS_01|0f|FL|1|Z tracking Error
0045|GEMS_HELIOS_01|10|SS|1|Start View 2A
0045|GEMS_HELIOS_01|11|SS|1|Number of Views 2A
0045|GEMS_HELIOS_01|12|SS|1|Start View 1A
0045|GEMS_HELIOS_01|13|SS|1|Sigma Mode
0045|GEMS_HELIOS_01|14|SS|1|Number of Views 1A
0045|GEMS_HELIOS_01|15|SS|1|Start View 2B
0045|GEMS_HELIOS_01|16|SS|1|Number Views 2B
0045|GEMS_HELIOS_01|17|SS|1|Start View 1B
0045|GEMS_HELIOS_01|21|SS|1|Iterbone Flag
0045|GEMS_HELIOS_01|22|SS|1|PeristalticFlag
0045|GEMS_HELIOS_01|30|CS|1|CardiacReconAlgorithm
0045|GEMS_HELIOS_01|31|CS|1|AvgHeartRateForImage
0045|GEMS_HELIOS_01|32|FL|1|TemporalResolution
0045|GEMS_HELIOS_01|33|CS|1|PctRpeakDelay
0045|GEMS_HELIOS_01|36|CS|1|EkgFullMaStartPhase
0045|GEMS_HELIOS_01|37|CS|1|EkgFullMaEndPhase
0045|GEMS_HELIOS_01|38|CS|1|EkgModulationMaxMa
0045|GEMS_HELIOS_01|39|CS|1|EkgModulationMinMa
0045|GEMS_HELIOS_01|3b|LO|1|NoiseReductionImageFilterDesc
0047|GEMS_IQTB_IDEN_47|02|UL|1|Unknown
0119|MRSC|1201|LO|1|SourceID
004b|GEMS_CT_HINO_01|01|DS|1-n|Beam Thickess
004b|GEMS_CT_HINO_01|02|DS|1-n|R Time
004b|GEMS_CT_HINO_01|03|IS|1|HBC Number
004b|GEIIS|13|IS|1|Unknown
004b|GEIIS|15|LT|1|Unknown
0051|GEMS_CT_VES_01|01|SQ|1|CTVESequence
0055|GEMS_GENIE_1|12|SQ|1|eNTEGRA Energy Window Information Sequence
0055|GEMS_GENIE_1|13|SQ|1|eNTEGRA Energy Window Range Sequence
0055|GEMS_GENIE_1|22|SQ|1|eNTEGRA Detector Information Sequence
0055|GEMS_GENIE_1|52|SQ|1|eNTEGRA Rotation Information Sequence
0055|GEMS_GENIE_1|62|SQ|1|eNTEGRA Gated Information Sequence
0055|GEMS_GENIE_1|63|SQ|1|eNTEGRA Data Information Sequence
0055|GEMS_GENIE_1|64|SQ|1|SDO Double Data Sequence
0055|GEMS_GENIE_1|65|SQ|1|Unknown
3101|AMI Annotations_01|10|SQ|1|Annotation Sequence
3101|AMI Annotations_02|20|SQ|1|Annotation Sequence
3103|AMI Sequence Annotations_01|10|CS|1|Annotation Sequence
3103|AMI Sequence Annotations_01|20|UI|1|Annotation UID
3103|AMI Sequence Annotations_01|30|US|1|Annotation Color
3103|AMI Sequence Annotations_01|50|CS|1|Annotation Line Style
3103|AMI Sequence Annotations_01|60|SQ|1|Annotation Elements
3103|AMI Sequence Annotations_01|70|SH|1|Annotation Label
3103|AMI Sequence Annotations_01|80|PN|1|Annotation Creator
3103|AMI Sequence Annotations_01|90|PN|1|Annotation Modifiers
3103|AMI Sequence Annotations_01|a0|DA|1|Annotation Creation Date
3103|AMI Sequence Annotations_01|b0|TM|1|Annotation Creation Time
3103|AMI Sequence Annotations_01|c0|DA|1|Annotation Modification Dates
3103|AMI Sequence Annotations_01|d0|TM|1|Annotation Mofification Times
3103|AMI Sequence Annotations_01|e0|US|1|Annotation Frame Number
3103|AMI Sequence Annotations_02|10|CS|1|Annotation Sequence
3103|AMI Sequence Annotations_02|20|UI|1|Annotation UID
3103|AMI Sequence Annotations_02|30|US|1|Annotation Color
3103|AMI Sequence Annotations_02|50|CS|1|Annotation Line Style
3103|AMI Sequence Annotations_02|60|SQ|1|Annotation Elements
3103|AMI Sequence Annotations_02|70|SH|1|Annotation Label
3103|AMI Sequence Annotations_02|80|PN|1|Annotation Creator
0049|GEMS_CT_CARDIAC_001|02|CS|1|HeartRateAtConfirm
0049|GEMS_CT_CARDIAC_001|03|FL|1|AvgHeartRatePriorToConfirm
0049|GEMS_CT_CARDIAC_001|04|CS|1|MinHeartRatePriorToConfirm
0049|GEMS_CT_CARDIAC_001|06|FL|1|StdDevHeartRatePriorToConfirm
0049|GEMS_CT_CARDIAC_001|07|US|1|NumHeartRateSamplesPriorToConfirm
0049|GEMS_CT_CARDIAC_001|08|CS|1|AutoHeartRateDetectPredict
0049|GEMS_CT_CARDIAC_001|09|CS|1|SystemOptimizedHeartRate
0049|GEMS_CT_CARDIAC_001|0a|ST|1|EkgMonitorType
0049|GEMS_CT_CARDIAC_001|0b|CS|1|NumReconSectors
0049|GEMS_CT_CARDIAC_001|0c|FL|256|RpeakTimeStamps
3103|AMI Sequence Annotations_02|90|PN|1|Annotation Modifiers
3103|AMI Sequence Annotations_02|a0|DA|1|Annotation Creation Date
3103|AMI Sequence Annotations_02|b0|TM|1|Annotation Creation Time
3103|AMI Sequence Annotations_02|c0|DA|1|Annotation Modification Dates
3103|AMI Sequence Annotations_02|d0|TM|1|Annotation Modification Times
3103|AMI Sequence Annotations_02|e0|US|1|Annotation Frame Number
3105|AMI Sequence AnnotElements_01|10|DS|1-n|Annotation Element Position
3105|AMI Sequence AnnotElements_01|20|LT|1|Annotation Element Text
3107|AMI ImageTransform_01|10|DS|1-n|Transformation Matrix
3107|AMI ImageTransform_01|20|DS|1|Center Offset
3107|AMI ImageTransform_01|30|DS|1|Magnification
3107|AMI ImageTransform_01|40|CS|1|Magnification Type
3107|AMI ImageTransform_01|50|DS|1|Displayed Area
3107|AMI ImageTransform_01|60|DS|1|Calibration Factor
3107|AMI ImageContextExt_01|a0|CS|1|Window Function
3107|AMI ImageContextExt_01|b0|DS|1|Window Slope
3109|Applicare/RadWorks/Version 5.0|01|ST|1|Worklist Filename
3109|Applicare/RadWorks/Version 5.0|02|SH|1|NEW/SEEN Status
3109|Applicare/RadWorks/Version 5.0|03|CS|1|Delete Lock
3109|Applicare/RadWorks/Version 5.0|04|CS|1|Unknown
3109|Applicare/RadWorks/Version 5.0|05|CS|1|Unknown
3109|Applicare/RadWorks/Version 5.0|06|CS|1|Unknown
3109|Applicare/RadWorks/Version 5.0|07|UL|1|Unknown
3109|Applicare/RadWorks/Version 5.0|08|LO|1|Receive Origin
3109|Applicare/RadWorks/Version 5.0|09|LO|1|Folder
3109|Applicare/RadWorks/Version 5.0|0a|DA|1|Receive Date
3109|Applicare/RadWorks/Version 5.0|0b|TM|1|Receive Time
3109|Applicare/RadWorks/Version 5.0|0c|CS|1|Prior
3109|Applicare/RadWorks/Version 5.0|0d|CS|1|STAT Study
3109|Applicare/RadWorks/Version 5.0|0e|CS|1|Is Key Image Or Study
3109|Applicare/RadWorks/Version 5.0|10|CS|1|Local Study
3109|Applicare/RadWorks/Version 5.0|11|LO|1|Result Message
3109|Applicare/RadWorks/Version 5.0|12|LO|1|Current User
3109|Applicare/RadWorks/Version 5.0|13|DA|1|System Date
3109|Applicare/RadWorks/Version 5.0|14|TM|1|System Time
3109|Applicare/RadWorks/Version 5.0|19|LO|1|Worklist Name
3109|Applicare/RadWorks/Version 5.0|20|UI|1|Worklist UID
3109|Applicare/RadWorks/Version 5.0|21|CS|1|Hostname
3109|Applicare/RadWorks/Version 5.0|22|AE|1|DICOM AE Title
3109|Applicare/RadWorks/Version 5.0|23|US|1|DICOM Port Number
3109|Applicare/RadWorks/Version 5.0|24|LO|1|Destination Name
3109|Applicare/RadWorks/Version 5.0|25|LO|1|Origin Name
3109|Applicare/RadWorks/Version 5.0|26|UI|1|Modality Study Instance UID
3109|Applicare/RadWorks/Version 5.0|27|SQ|1|Exam Routing
3109|Applicare/RadWorks/Version 5.0|28|LO|1|Notification Comments
3109|Applicare/RadWorks/Version 5.0|29|LO|1|Transaction Comments
3109|Applicare/RadWorks/Version 5.0|2a|LO|1|Send Flag
3109|Applicare/RadWorks/Version 5.0|2b|LO|1|Print Flag
3109|Applicare/RadWorks/Version 5.0|2c|LO|1|Archive Flag
3109|Applicare/RadWorks/Version 5.0|30|LO|1|Requesting Facility Name
3109|Applicare/RadWorks/Version 5.0|31|CS|1|Requesting Procedure Name
3109|Applicare/RadWorks/Version 5.0|32|CS|1|Requesting Procedure Code
3109|Applicare/RadWorks/Version 5.0|33|CS|1|Request Storage Commitment
3109|Applicare/RadWorks/Version 5.0|34|CS|1|Requested Compression
3109|Applicare/RadWorks/Version 5.0|35|SQ|1|Study Sequence
3109|Applicare/RadWorks/Version 5.0|37|UI|1|Replaced Study UID
3109|Applicare/RadWorks/Version 5.0|38|SH|1|Teaching ACR Code
3109|Applicare/RadWorks/Version 5.0|39|SH|1|Teaching Special Interest Code
3109|Applicare/RadWorks/Version 5.0|40|IS|1|Number of Study Related Images
3109|Applicare/RadWorks/Version 5.0|41|CS|1|Study Locked
3109|Applicare/RadWorks/Version 5.0|42|CS|1|Workstation Name
3109|Applicare/RadWorks/Version 5.0|43|CS|1|Archive Status
3109|Applicare/RadWorks/Version 5.0|ee|UI|1|Internal List UID
3109|Applicare/RadWorks/Version 5.0|ef|CS|1|Action (Add,Remove,Change)
3109|Applicare/RadWorks/Version 6.0/Summary|01|SH|1|Status
3109|Applicare/RadWorks/Version 6.0/Summary|11|ST|1|Receive Origin Site Name
3109|Applicare/RadWorks/Version 6.0/Summary|12|ST|1|Receive Origin Description
3109|Applicare/RadWorks/Version 6.0/Summary|15|DA|1|Receive Date
3109|Applicare/RadWorks/Version 6.0/Summary|16|TM|1|Receive Time
3115|http://www.gemedicalsystems.com/it_solutions/rad_pacs/|01|UT|1|Unknown
4101|Applicare/Print/Version 5.1|01|UL|1|Mask State
4101|Applicare/Print/Version 5.1|02|SQ|1|Annotations
4101|Applicare/Print/Version 5.1|03|LO|1|Font
4101|Applicare/Print/Version 5.1|04|UL|1|Font Size
4101|Applicare/Print/Version 5.1|05|FD|1|Font Relative Size
4101|Applicare/Print/Version 5.1|06|US|1|Overlay
4101|Applicare/Print/Version 5.1|07|US|1|Pixel Rep
4101|Applicare/Print/Version 5.1|08|US|1|Annotation Level
4101|Applicare/Print/Version 5.1|09|US|1|Show Caliper
4103|Applicare/RadWorks/Version 6.0|01|AT|1-n|Non-existent tags
4103|Applicare/RadWorks/Version 6.0|02|UI|1-n|Non-existent objects
4105|Applicare/RadWorks/Version 6.0|01|CS|1|Annotation Type
4105|Applicare/RadWorks/Version 6.0|02|LO|1|Annotation Value
4105|Applicare/RadWorks/Version 6.0|03|UI|1|Cutline Image UID
4105|Applicare/RadWorks/Version 6.0|04|UI|1|Cutline Set UID
5001|GEMS_GENIE_1|35|LO|1|Dataset Name
4105|Applicare/RadWorks/Version 6.0|05|US|3|Annotation Color (RGB)
4105|Applicare/RadWorks/Version 6.0|06|CS|1|Annotation Line Style
4105|Applicare/RadWorks/Version 6.0|07|SH|1|Annotation Label
4105|Applicare/RadWorks/Version 6.0|08|PN|1|Annotation Creator
4105|Applicare/RadWorks/Version 6.0|09|DA|1|Annotation Creation Date
4105|Applicare/RadWorks/Version 6.0|0a|TM|1|Annotation Creation Time
4105|Applicare/RadWorks/Version 6.0|0b|SQ|1|Annotation Modification Sequence
4105|Applicare/RadWorks/Version 6.0|0c|PN|1|Annotation Modifier
4105|Applicare/RadWorks/Version 6.0|0d|DA|1|Annotation Modification Date
4105|Applicare/RadWorks/Version 6.0|0e|TM|1|Annotation Modification Time
4105|Applicare/RadWorks/Version 6.0|10|US|1|Unknown
4107|Applicare/RadWorks/Version 6.0|01|SQ|1|Requested Palette Color LUT
5001|GEMS_GENIE_1|01|SL|1|Modified
5001|GEMS_GENIE_1|02|LO|1|Name
5001|GEMS_GENIE_1|03|SL|1|Cid
5001|GEMS_GENIE_1|04|SL|1|Srid
5001|GEMS_GENIE_1|05|LO|1|SOP Class UID
5001|GEMS_GENIE_1|06|LO|1|SOP Instance UID
5001|GEMS_GENIE_1|07|SL|1|Curve Type
5001|GEMS_GENIE_1|08|SL|1|Graph Type
5001|GEMS_GENIE_1|09|LO|1|Legend
5001|GEMS_GENIE_1|0a|LO|1|X Units
5001|GEMS_GENIE_1|0b|LO|1|Y Units
5001|GEMS_GENIE_1|0c|SL|1|Edit
5001|GEMS_GENIE_1|0d|SL|1|Suspend
5001|GEMS_GENIE_1|0e|SL|1|Style Line
5001|GEMS_GENIE_1|0f|SL|1|Style Fill
5001|GEMS_GENIE_1|10|LO|1|Style Colour
5001|GEMS_GENIE_1|11|SL|1|Style Width
5001|GEMS_GENIE_1|12|SL|1|Style Point
5001|GEMS_GENIE_1|13|LO|1|Style P Colour
5001|GEMS_GENIE_1|14|SL|1|Style P Size
5001|GEMS_GENIE_1|15|SL|1|Segments
5001|GEMS_GENIE_1|16|SL|1|Seg Type
5001|GEMS_GENIE_1|17|FD|1-n|Seg Start
5001|GEMS_GENIE_1|18|FD|1-n|Seg End
5001|GEMS_GENIE_1|19|SL|1-n|Seg Style Line
5001|GEMS_GENIE_1|1a|SL|1-n|SegStyleFill
5001|GEMS_GENIE_1|1b|LO|1|Seg Style Colour
5001|GEMS_GENIE_1|1c|SL|1-n|Seg Style Width
5001|GEMS_GENIE_1|1d|SL|1-n|Seg Style Point
5001|GEMS_GENIE_1|1e|SL|1|Seg Style P Colour
5001|GEMS_GENIE_1|1f|SL|1|Seg Style P Size
5001|GEMS_GENIE_1|20|LO|1|Seg Name
5001|GEMS_GENIE_1|21|SL|1-n|Seg Allow Dir Int
5001|GEMS_GENIE_1|22|SL|1|Text Annots
5001|GEMS_GENIE_1|23|FD|1-n|Txt X
5001|GEMS_GENIE_1|24|FD|1-n|Txt Y
5001|GEMS_GENIE_1|25|LO|1|Txt Text
5001|GEMS_GENIE_1|26|LO|1|Txt Name
5001|GEMS_GENIE_1|30|LO|1|ROI Name
5001|GEMS_GENIE_1|31|LO|1|Derived From Image UID
5001|GEMS_GENIE_1|32|SL|1-n|Derived From Images
5001|GEMS_GENIE_1|33|UL|1|Curve Flags
5001|GEMS_GENIE_1|34|LO|1|Curve Name
5001|GEMS_GENIE_1|36|LO|1|Curve UID
5001|GEMS_GENIE_1|37|FD|1|ROI Area
5001|GEMS_GENIE_1|38|LO|1|Modified
5001|GEMS_GENIE_1|39|LO|1|Name
5001|GEMS_GENIE_1|3a|LO|1|Software Version
5001|GEMS_GENIE_1|3b|SH|1|Start Date
5001|GEMS_GENIE_1|3c|SH|1|Completion Date
5001|GEMS_GENIE_1|3d|LO|1|Detector Name
5001|GEMS_GENIE_1|41|SL|1|Modified
5001|GEMS_GENIE_1|42|LO|1|Name
5001|GEMS_GENIE_1|43|SL|1|Name
5001|GEMS_GENIE_1|44|SL|1|Name
5001|GEMS_GENIE_1|45|LO|1|SOP Class UID
5001|GEMS_GENIE_1|46|LO|1|SOP Instance UID
5001|GEMS_GENIE_1|47|LO|1|Normal Color
5001|GEMS_GENIE_1|48|LT|1|Name Font
5001|GEMS_GENIE_1|49|SL|1|Fill Pattern
5001|GEMS_GENIE_1|4a|SL|1|Line Style
5001|GEMS_GENIE_1|4b|SL|1|Line Dash Length
5001|GEMS_GENIE_1|4c|SL|1|Line Thickness
5001|GEMS_GENIE_1|4d|SL|1|Interactivity
5001|GEMS_GENIE_1|4e|SL|1|Name Pos
5001|GEMS_GENIE_1|4f|SL|1|Name Display
5001|GEMS_GENIE_1|50|LO|1|Label
5001|GEMS_GENIE_1|51|SL|1-n|Bp Seg
5001|GEMS_GENIE_1|52|US|1-n|Bp Seg Pairs
5001|GEMS_GENIE_1|53|SL|1|Seed Space
5001|GEMS_GENIE_1|54|FD|1-n|Seeds
5001|GEMS_GENIE_1|55|SL|1-n|Shape
5001|GEMS_GENIE_1|56|FD|1-n|Shape Tilt
5001|GEMS_GENIE_1|59|SL|1-n|Shape Pts Space
5001|GEMS_GENIE_1|5a|SL|1-n|Shape Ctrl Pts Counts
5001|GEMS_GENIE_1|5b|FD|1-n|Shape Ctrl Pts
5001|GEMS_GENIE_1|5c|SL|1|Shape Ctrl P Space
5001|GEMS_GENIE_1|5d|SL|1|ROI Flags
5001|GEMS_GENIE_1|5e|SL|1|Frame Number
5001|GEMS_GENIE_1|5f|SL|1|ID
5001|GEMS_GENIE_1|60|LO|1-n|Dataset ROI Mapping
0009|GEIIS|10|SQ|1|GE Private Image Thumbnail Sequence
0009|GEIIS|12|IS|1|Unknown
0029|GEIIS|10|UL|1|Shift Count
0029|GEIIS|12|UL|1|Offset
0029|GEIIS|14|UL|1|Actual Frame Number
0903|GEIIS PACS|10|US|1|Reject Image Flag
0903|GEIIS PACS|11|US|1|Significant Flag
0903|GEIIS PACS|12|US|1|Confidential Flag
0903|GEIIS PACS|20|CS|1|Unknown
0905|GEIIS|30|LO|1|Assigning Authority For Patient ID
0907|GEIIS|10|UI|1|Original Study Instance UID
0907|GEIIS|20|UI|1|Original Series Instance UID
0907|GEIIS PACS|21|US|1|Prefetch Algorithm
0907|GEIIS PACS|22|US|1|Limit Recent Studies
0907|GEIIS PACS|23|US|1|Limit Oldest Studies
0907|GEIIS PACS|24|US|1|Limit Recent Months
0907|GEIIS|30|UI|1|Original SOP Instance UID
0907|GEIIS PACS|31|UI|1-n|Exclude Study UIDs
7fd1|GEIIS|10|UL|1|Compression Type
7fd1|GEIIS|20|UL|1-n|Multiframe Offsets
7fd1|GEIIS|30|UL|1|Multi-Resolution Levels
7fd1|GEIIS|40|UL|1-n|Subband Rows
7fd1|GEIIS|50|UL|1-n|Subband Columns
7fd1|GEIIS|60|UL|1-n|Subband Bytecounts
0011|GEMS_GDXE_FALCON_04|03|UI|1|Processed Series UID
0011|GEMS_GDXE_FALCON_04|04|CS|1|Acquisition Type
0011|GEMS_GDXE_FALCON_04|05|UI|1|Acquisition UID
0011|GEMS_GDXE_FALCON_04|06|DS|1|Image Dose
0011|GEMS_GDXE_FALCON_04|07|FL|1|Study Dose
0011|GEMS_GDXE_FALCON_04|08|FL|1|Study DAP
0011|GEMS_GDXE_FALCON_04|09|SL|1|Non-Digital Exposures
0011|GEMS_GDXE_FALCON_04|10|SL|1|Total Exposures
0011|GEMS_GDXE_FALCON_04|11|LT|1|ROI
0011|GEMS_GDXE_FALCON_04|12|LT|1|Patient Size String
0011|GEMS_GDXE_FALCON_04|13|UI|1|SPS UID
0011|GEMS_GDXE_FALCON_04|14|UI|1|Unknown
0011|GEMS_GDXE_FALCON_04|15|DS|1|Detector ARC Gain
0011|GEMS_GDXE_FALCON_04|16|LT|1|Processing Debug Info
0011|GEMS_GDXE_FALCON_04|17|CS|1|Override Mode
0011|GEMS_GDXE_FALCON_04|19|DS|1|Film Speed Selection
0011|GEMS_GDXE_FALCON_04|27|UN|1|Unknown
0011|GEMS_GDXE_FALCON_04|28|UN|1|Unknown
0011|GEMS_GDXE_FALCON_04|29|UN|1|Unknown
0011|GEMS_GDXE_FALCON_04|30|UN|1|Unknown
0011|GEMS_GDXE_FALCON_04|31|IS|1-n|Detected Field of View
0011|GEMS_GDXE_FALCON_04|32|IS|1-n|Adjusted Field of View
0011|GEMS_GDXE_FALCON_04|33|DS|1|Detector Exposure Index
0011|GEMS_GDXE_FALCON_04|34|DS|1|Compensated Detector Exposure
0011|GEMS_GDXE_FALCON_04|35|DS|1|Uncompensated Detector Exposure
0011|GEMS_GDXE_FALCON_04|36|DS|1|Median Anatomy Count Value
0011|GEMS_GDXE_FALCON_04|37|DS|2|DEI Lower & Upper Limit Values
0011|GEMS_GDXE_FALCON_04|38|SL|6|Shift Vector for Pasting
0011|GEMS_GDXE_FALCON_04|39|CS|6|Image Number in Pasting
0011|GEMS_GDXE_FALCON_04|40|SL|1|Pasting Overlap
0011|GEMS_GDXE_FALCON_04|41|IS|24|Sub-image Collimator Vertices
0011|GEMS_GDXE_FALCON_04|42|LO|1|View IP
0011|GEMS_GDXE_FALCON_04|43|IS|24|Keystone Coordinates
0011|GEMS_GDXE_FALCON_04|44|CS|1|Receptor Type
0011|GEMS_GDXE_FALCON_04|46|LO|1-n|Unknown
0011|GEMS_GDXE_FALCON_04|47|DS|1|Unknown
0011|GEMS_GDXE_FALCON_04|59|CS|1|Unknown
0011|GEMS_GDXE_FALCON_04|60|CS|1|Unknown
0011|GEMS_GDXE_FALCON_04|6d|DS|1|Unknown
0045|GEMS_FALCON_03|55|DS|8|A_Coefficients used in Multiresolution Algorithm
0045|GEMS_FALCON_03|62|IS|1|User Window Center
0045|GEMS_FALCON_03|63|IS|1|User Window Width
0045|GEMS_FALCON_03|65|IS|1|Requested Detector Entrance Dose
0045|GEMS_FALCON_03|67|DS|3|VOI LUT Assymmetry Parameter Beta
0045|GEMS_FALCON_03|69|IS|1|Collimator Rotation
0045|GEMS_FALCON_03|72|IS|1|Collimator Width
0045|GEMS_FALCON_03|73|IS|1|Collimator Height
0045|GEMS_SEND_02|55|DS|8|A_Coefficients used in Multiresolution Algorithm
0045|GEMS_SEND_02|62|IS|1|User Window Center
0045|GEMS_SEND_02|63|IS|1|User Window Width
0045|GEMS_SEND_02|65|IS|1|Requested Detector Entrance Dose
0045|GEMS_SEND_02|67|DS|3|VOI LUT Assymmetry Parameter Beta
0045|GEMS_SEND_02|69|IS|1|Collimator Rotation
0045|GEMS_SEND_02|72|IS|1|Collimator Width
0045|GEMS_SEND_02|73|IS|1|Collimator Height
7fdf|GEMS_GDXE_ATHENAV2_INTERNAL_USE|10|LT|1|Pixel Data References
7fdf|GEMS_GDXE_ATHENAV2_INTERNAL_USE|11|LT|1|Pixel Data References (temporary)
7fdf|GEMS_GDXE_ATHENAV2_INTERNAL_USE|20|SS|1|Auto Push Tag
7fdf|GEMS_GDXE_ATHENAV2_INTERNAL_USE|25|CS|1|PPS Status
6003|GEMS_Ultrasound_ImageGroup_001|10|SQ|1|Unknown
6003|GEMS_Ultrasound_ImageGroup_001|11|OB|1|Unknown
6003|GEMS_Ultrasound_ImageGroup_001|12|LT|1|Unknown
6003|GEMS_Ultrasound_ImageGroup_001|15|LT|1-n|Unknown
6005|GEMS_Ultrasound_ExamGroup_001|10|UT|1|Unknown
6005|GEMS_Ultrasound_ExamGroup_001|20|UT|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|01|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|02|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|03|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|08|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|10|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|12|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|18|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|20|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|24|SH|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|26|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|30|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|32|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|36|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|37|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|3a|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|3c|FD|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|43|OB|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|48|FD|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|49|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|51|FL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|52|FD|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|53|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|54|SL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|55|OB|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|57|LT|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|60|OB|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|61|OW|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|62|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|69|OW|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|70|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|71|UL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|72|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|73|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|74|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|75|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|77|FD|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|79|SL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|83|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|84|LO|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|85|SQ|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|86|SL|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|87|FD|1|Unknown
7fe1|GEMS_Ultrasound_MovieGroup_001|88|FD|1|Unknown
7fe1|KRETZ_US|01|OB|1|Unknown
0009|QUASAR_INTERNAL_USE|01|UL|1-n|Rate Vector
0009|QUASAR_INTERNAL_USE|02|UL|1-n|Count Vector
0009|QUASAR_INTERNAL_USE|03|UL|1-n|Time Vector
0009|QUASAR_INTERNAL_USE|07|UL|1-n|Angle Vector
0009|QUASAR_INTERNAL_USE|08|US|1|Camera Shape
0009|QUASAR_INTERNAL_USE|10|US|1|Whole Body Spots
0009|QUASAR_INTERNAL_USE|11|US|1|Worklist Flag
0009|QUASAR_INTERNAL_USE|12|LO|1|Unknown
0009|QUASAR_INTERNAL_USE|13|ST|1|Sequence Type
0009|QUASAR_INTERNAL_USE|14|ST|1|Sequence Name
0009|QUASAR_INTERNAL_USE|15|UL|1-n|Average RR Time Vector
0009|QUASAR_INTERNAL_USE|16|UL|1-n|Low Limit Vector
0009|QUASAR_INTERNAL_USE|17|UL|1-n|High Limit Vector
0009|QUASAR_INTERNAL_USE|18|UL|1-n|Begin Index Vector
0009|QUASAR_INTERNAL_USE|19|UL|1-n|End Index Vector
0009|QUASAR_INTERNAL_USE|1a|UL|1-n|Raw Time Vector
0009|QUASAR_INTERNAL_USE|1b|LO|1|Image Type String
0009|QUASAR_INTERNAL_USE|1d|US|1|Unknown
0009|QUASAR_INTERNAL_USE|1e|ST|1|Unknown
0009|QUASAR_INTERNAL_USE|22|FL|1|Unknown
0009|QUASAR_INTERNAL_USE|23|US|1|Unknown
0009|QUASAR_INTERNAL_USE|39|UI|1|Unknown
0009|QUASAR_INTERNAL_USE|40|DA|1|Unknown
0009|QUASAR_INTERNAL_USE|41|TM|1|Unknown
0009|QUASAR_INTERNAL_USE|42|LO|1|Unknown
0009|QUASAR_INTERNAL_USE|44|SH|1|Unknown
0009|QUASAR_INTERNAL_USE|45|LO|1|Unknown
0009|QUASAR_INTERNAL_USE|48|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|10|SQ|1|Unknown
0037|QUASAR_INTERNAL_USE|1b|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|30|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|40|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|50|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|60|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|70|LO|1|Unknown
0037|QUASAR_INTERNAL_USE|71|FD|1|Unknown
0037|QUASAR_INTERNAL_USE|72|SH|1|Unknown
0037|QUASAR_INTERNAL_USE|73|FD|1|Unknown
0037|QUASAR_INTERNAL_USE|78|FD|1|Unknown
0037|QUASAR_INTERNAL_USE|90|IS|1|Unknown
0037|QUASAR_INTERNAL_USE|92|DS|1|Unknown
0041|QUASAR_INTERNAL_USE|01|UT|1|Unknown
0027|APEX_PRIVATE|11|DS|1|Bed Position
0033|GEMS_XELPRV_01|08|CS|1|Unknown
0033|GEMS_XELPRV_01|10|SL|1|Unknown
0033|GEMS_XELPRV_01|11|LO|1|Unknown
0033|GEMS_XELPRV_01|16|UI|1|Unknown
0033|GEMS_XELPRV_01|17|DA|1|Unknown
0033|GEMS_XELPRV_01|18|TM|1|Unknown
0033|GEMS_XELPRV_01|19|UL|1|Unknown
0033|GEMS_XELPRV_01|1a|LO|1|Unknown
0033|GEMS_XELPRV_01|1b|LO|1|Unknown
0033|GEMS_XELPRV_01|1c|OB|1|Unknown
0033|GEMS_XELPRV_01|1d|UL|1|Unknown
0033|GEMS_XELPRV_01|1e|FD|1|Unknown
0033|GEMS_XELPRV_01|1f|OB|1|Unknown
0033|GEMS_XELPRV_01|20|OB|1|Unknown
0033|GEMS_XELPRV_01|21|OB|1|Unknown
0033|GEMS_XELPRV_01|22|OB|1|Unknown
0033|GEMS_XELPRV_01|23|OB|1|Unknown
0033|GEMS_XELPRV_01|24|LT|1|Unknown
0033|GEMS_XELPRV_01|70|SQ|1|Unknown
0033|GEMS_XELPRV_01|71|UI|1|Unknown
0033|GEMS_XELPRV_01|72|UI|1|Unknown
0039|REPORT_FROM_APP|95|LO|1|Unknown
0047|GEMS_VXTL_USERDATA_01|11|LT|1|Unknown
0015|DL_INTERNAL_USE|8f|IS|1|Unknown
7003|GEMS_LUNAR_RAW|01|ST|1|enCORE File Name
7003|GEMS_LUNAR_RAW|02|OB|1|enCORE File Data
7003|GEMS_LUNAR_RAW|03|UL|1|enCORE File Length
7003|GEMS_LUNAR_RAW|04|LO|1|enCORE File Modified Time
0119|MRSC|1202|IS|1|Group Version
6005|GE_GROUP|10|UT|1|Unknown
0087|1.2.840.113708.794.1.1.2.0|30|ST|1|Storage File ID
0087|1.2.840.113708.794.1.1.2.0|40|DS|1|Study or Image Size in MB
0045|GEMS_IT_US_REPORT|11|OW|1|Vivid excel file
0045|GEMS_IT_US_REPORT|12|OW|1|Vivid CHM file
0045|GEMS_IT_US_REPORT|13|OW|1|Vivid PDF file
3113|Applicare/Workflow/Version 1.0|01|CS|1|Order Control
3113|Applicare/Workflow/Version 1.0|10|SH|1|Scheduled Action Item Code Value
3113|Applicare/Workflow/Version 1.0|11|SH|1|Scheduled Action Item Coding Scheme Designator
3113|Applicare/Workflow/Version 1.0|12|LO|1|Scheduled Action Item Code Meaning
3113|Applicare/Workflow/Version 1.0|15|SH|1|Requested Action Item Code Value
3113|Applicare/Workflow/Version 1.0|16|SH|1|Requested Action Item Coding Scheme Designator
0053|GEHC_CT_ADVAPP_001|20|IS|1|Shuttle Flag
0053|GEHC_CT_ADVAPP_001|40|SH|1|Iterative Recon Annotation
0053|GEHC_CT_ADVAPP_001|41|SH|1|Iterative Recon Mode
0053|GEHC_CT_ADVAPP_001|42|LO|1|Iterative Recon Configuration
0053|GEHC_CT_ADVAPP_001|43|SH|1|Iterative Recon Level
0053|GEHC_CT_ADVAPP_001|61|SH|1|High Resolution Flag
0053|GEHC_CT_ADVAPP_001|62|SH|1|Respiratory Flag
0053|GEHC_CT_ADVAPP_001|9d|LO|1|Unknown
3113|Applicare/Workflow/Version 1.0|17|LO|1|Requested Action Item Code Meaning
3113|Applicare/Workflow/Version 1.0|20|SH|1|Performed Action Item Code Value
3113|Applicare/Workflow/Version 1.0|21|SH|1|Performed Action Item Coding Scheme Designator
3113|Applicare/Workflow/Version 1.0|22|LO|1|Performed Action Item Code Meaning
3113|Applicare/Workflow/Version 1.0|25|SH|1|Performed Procedure Code Value
3113|Applicare/Workflow/Version 1.0|26|SH|1|Performed Procedure Coding Scheme Designator
3113|Applicare/Workflow/Version 1.0|27|LO|1|Performed Procedure Code Meaning
3113|Applicare/Workflow/Version 1.0|30|UI|1|Referenced Image SOP Class UID
3113|Applicare/Workflow/Version 1.0|31|UI|1|Referenced Image SOP Instance UID
3113|Applicare/Workflow/Version 1.0|e0|CS|1|Locked By Hostname
3113|Applicare/Workflow/Version 1.0|e1|CS|1|Locked By User
3113|Applicare/Workflow/Version 1.0|e2|CS|1|KfEdit Lock User
0045|GE LUT Asymmetry Parameter|67|DS|1|LUT Assymetry
4109|Applicare/Centricity Radiology Web/Version 1.0|01|SH|1|Mammography Laterality
4109|Applicare/Centricity Radiology Web/Version 1.0|02|SH|1|Mammography View Name
4109|Applicare/Centricity Radiology Web/Version 1.0|03|SH|1|Mammography View Modifier
4111|Applicare/Centricity Radiology Web/Version 2.0|01|CS|1|Secondary Spine Label
4111|Applicare/Centricity Radiology Web/Version 2.0|02|IS|1|Additional tags for Presentation State
4113|GEMS-IT/Centricity RA600/7.0|10|UI|1|Number of images in study
3111|AMI StudyExtensions_01|01|UL|1|Last Released Annot Label
3111|RadWorksTBR|02|CS|1|Compression Type
3111|RadWorksTBR|ff|SQ|1|Query Result
3113|Applicare/RadStore/Version 1.0|01|SL|1|Unknown
3113|Applicare/RadStore/Version 1.0|02|SL|1|Internal Id of Study
3113|Applicare/RadStore/Version 1.0|03|SL|1|Internal Id of Series
3113|Applicare/RadStore/Version 1.0|04|SL|1|Internal Id of Instance
3113|Applicare/RadStore/Version 1.0|11|LO|1|Unknown
3113|Applicare/RadStore/Version 1.0|12|CS|1|Instance State
3113|Applicare/RadStore/Version 1.0|13|DT|1|Date Last Modified
3113|Applicare/RadStore/Version 1.0|14|DT|1|Date Last Accessed
3113|Applicare/RadStore/Version 1.0|15|CS|1|Unknown
3113|Applicare/RadStore/Version 1.0|16|FD|1|Instance Size in Bytes
3113|Applicare/RadStore/Version 1.0|17|LO|1|Library Id
3113|Applicare/RadStore/Version 1.0|18|LO|1|Pathnames
3113|Applicare/RadStore/Version 1.0|19|LO|1|Driver Path
3113|Applicare/RadStore/Version 1.0|1a|LO|1|Source
3113|Applicare/RadStore/Version 1.0|1b|LO|1|Destination
3113|Applicare/RadStore/Version 1.0|1c|SL|1|Medium Id
3113|Applicare/RadStore/Version 1.0|1d|LO|1|Archive Id
3113|Applicare/RadStore/Version 1.0|1e|LO|1|Instance Origin
3113|Applicare/RadStore/Version 1.0|21|SL|1|Instance Version
3113|Applicare/RadStore/Version 1.0|22|SL|1|Unknown
3113|Applicare/RadStore/Version 1.0|23|ST|1|Instance File Location
3113|Applicare/RadStore/Version 1.0|31|IS|1|Unknown
3113|Applicare/RadStore/Version 1.0|32|IS|1|Unknown
3113|Applicare/RadStore/Version 1.0|33|IS|1|Unknown
3113|Applicare/RadStore/Version 1.0|35|LO|1|Image Medium Location
3113|Applicare/RadStore/Version 1.0|36|LO|1|Image Medium Label
3113|Applicare/RadStore/Version 1.0|37|CS|1|Image Medium State
3113|Applicare/RadStore/Version 1.0|38|LO|1|Series Medium Location
3113|Applicare/RadStore/Version 1.0|39|LO|1|Series Medium Label
3113|Applicare/RadStore/Version 1.0|3a|CS|1|Series Medium State
3113|Applicare/RadStore/Version 1.0|3b|LO|1|Study Medium Location
3113|Applicare/RadStore/Version 1.0|3c|LO|1|Study Medium Label
3113|Applicare/RadStore/Version 1.0|3d|CS|1|Study Medium State
3113|Applicare/RadStore/Version 1.0|52|CS|1|Study State
3113|Applicare/RadStore/Version 1.0|53|CS|1|Series State
3113|Applicare/RadStore/Version 1.0|55|CS|1|Image State Text
3113|Applicare/RadStore/Version 1.0|56|CS|1|Series State Text
3113|Applicare/RadStore/Version 1.0|57|CS|1|Study State Text
3113|Applicare/RadStore/Version 1.0|60|DT|1|Expiration
3113|Applicare/RadStore/Version 1.0|69|AT|1-n|Deleted Tags
3115|http://www.gemedicalsystems.com/it_solutions/rad_pacs/|02|UT|1|Reference to pacs image
3115|http://www.gemedicalsystems.com/it_solutions/rad_pacs/|03|CS|1|Pacs examnotes flag
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|10|DT|1|OrthoView Session Date/Time
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|20|PN|1|OrthoView Session Creator
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|30|CS|1|OrthoView Session Completion Flag
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|40|SQ|1|OrthoView File Sequence
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|50|ST|1|OrthoView File Name
3117|http://www.gemedicalsystems.com/it_solutions/orthoview/2.1|60|OB|1|OrthoView File Content
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|10|DT|1|BAM WallThickness Session Date/Time
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|20|PN|1|BAM WallThickness Session Creator
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|30|CS|1|BAM WallThickness Session Completion Flag
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|40|SQ|1|BAM WallThickness File Sequence
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|50|ST|1|BAM WallThickness File Name
3118|http://www.gemedicalsystems.com/it_solutions/bamwallthickness/1.0|60|OB|1|BAM WallThickness File Content
3109|AMI ImageContext_01|10|CS|1|Window Invert
3109|AMI ImageContext_01|20|IS|1|Window Center
3109|AMI ImageContext_01|30|IS|1|Window Width
3109|AMI ImageContext_01|40|CS|1|Pixel Aspect Ratio Swap
3109|AMI ImageContext_01|50|CS|1|Enable Averaging
3109|AMI ImageContext_01|60|CS|1|Quality
3109|AMI ImageContext_01|70|CS|1|Viewport Annotation Level
3109|AMI ImageContext_01|80|CS|1|Show Image Annotation
3109|AMI ImageContext_01|90|CS|1|Show Image Overlay
0119|MRSC|1203|IS|1|ExecuteOnRead
0051|GEMS_FUNCTOOL_01|0d|OB|1|Wizard State
0019|Harmony R1.0|00|IS|1|Unknown
0019|Harmony R1.0|01|LO|1|Unknown
0019|Harmony R1.0|02|US|1|Unknown
0019|Harmony R1.0|03|IS|1|Unknown
0019|Harmony R1.0|04|UN|1|Unknown
0019|Harmony R1.0|05|UN|1|Unknown
0019|Harmony R1.0|06|UN|1|Unknown
0019|Harmony R1.0|07|UN|1|Unknown
0019|Harmony R1.0|08|UN|1|Unknown
0019|Harmony R1.0|09|US|1|Unknown
0019|Harmony R1.0|0a|US|1|Unknown
0019|Harmony R1.0|0b|US|1|Unknown
0019|Harmony R1.0|0c|UN|1|Unknown
0019|Harmony R1.0|0d|UN|1|Unknown
0019|Harmony R1.0|0e|US|1|Unknown
0019|Harmony R1.0|0f|UN|1|Unknown
0019|Harmony R1.0|10|UN|1|Unknown
0019|Harmony R1.0|11|UN|1|Unknown
0019|Harmony R1.0|12|TM|1|Unknown
0019|Harmony R1.0|13|UN|1|Unknown
0019|Harmony R1.0|14|UN|1|Unknown
0019|Harmony R1.0|15|UN|1|Unknown
0019|Harmony R1.0|16|IS|1-n|Unknown
0019|Harmony R1.0|17|US|1|Unknown
0019|Harmony R1.0|18|UN|1|Unknown
0019|Harmony R1.0|19|US|1|Unknown
0019|Harmony R1.0|1a|US|1|Unknown
0019|Harmony R1.0|1b|US|1|Unknown
0019|Harmony R1.0|1c|US|1|Unknown
0019|Harmony R1.0|1d|IS|1|Unknown
0019|Harmony R1.0|1e|US|1|Unknown
0019|Harmony R1.0|1f|US|1|Unknown
0019|Harmony R1.0|20|US|1|Unknown
0019|Harmony R1.0|24|UN|1|Unknown
0019|Harmony R1.0|25|IS|1|Unknown
0019|Harmony R1.0|26|IS|1|Unknown
0019|Harmony R1.0|29|UN|1|Unknown
0019|Harmony R1.0|2a|US|1|Unknown
0019|Harmony R1.0|2b|UN|1|Unknown
0051|GEMS_FUNCTOOL_01|02|LO|1|Function Name
0051|GEMS_FUNCTOOL_01|03|SL|1|Bias
0051|GEMS_FUNCTOOL_01|04|FL|1|Scale
0051|GEMS_FUNCTOOL_01|05|SL|1|Parameter Count
0051|GEMS_FUNCTOOL_01|06|LT|1|Parameters
0051|GEMS_FUNCTOOL_01|07|LO|1|Version
0051|GEMS_FUNCTOOL_01|09|SL|1|Window Width
0051|GEMS_FUNCTOOL_01|0a|SL|1|Window Level
0051|GEMS_FUNCTOOL_01|0b|FL|1|B-Value
0051|GEMS_FUNCTOOL_01|0c|SL|1|Wizard State Data Size
0019|Harmony R1.0|2d|UN|1|Unknown
0019|Harmony R1.0|2e|UN|1|Unknown
0019|Harmony R1.0|2f|UN|1|Unknown
0019|Harmony R1.0|30|UN|1|Unknown
0019|Harmony R1.0|31|UN|1|Unknown
0019|Harmony R1.0|32|UN|1|Unknown
0019|Harmony R1.0|33|UN|1|Unknown
0019|Harmony R1.0|34|UN|1|Unknown
0019|Harmony R1.0|35|UN|1|Unknown
0019|Harmony R1.0|36|UN|1|Unknown
0019|Harmony R1.0|37|UN|1|Unknown
0019|Harmony R1.0|38|UN|1|Unknown
0019|Harmony R1.0|39|UN|1|Unknown
0019|Harmony R1.0|3a|UN|1|Unknown
0019|Harmony R1.0|3b|US|1|Unknown
0019|Harmony R1.0|3c|US|1|Unknown
0019|Harmony R1.0|3d|UN|1|Unknown
0019|Harmony R1.0|3e|US|1|Unknown
0019|Harmony R1.0|3f|US|1|Unknown
0019|Harmony R1.0|40|UN|1|Unknown
0019|Harmony R1.0|41|UN|1|Unknown
0019|Harmony R1.0|42|LO|1|Unknown
0019|Harmony R1.0|43|US|1|Unknown
0019|Harmony R1.0|44|US|1|Unknown
0019|Harmony R1.0|45|UN|1|Unknown
0019|Harmony R1.0|46|US|1|Unknown
0019|Harmony R1.0|47|LO|1|Unknown
0019|Harmony R1.0|48|US|1|Unknown
0019|Harmony R1.0|49|US|1|Unknown
0019|Harmony R1.0|4a|US|1|Unknown
0019|Harmony R1.0|4b|UN|1|Unknown
0019|Harmony R1.0|4c|UN|1|Unknown
0019|Harmony R1.0|4e|UN|1|Unknown
0019|Harmony R1.0|4f|UN|1|Unknown
0019|Harmony R1.0|50|US|1|Unknown
0019|Harmony R1.0|51|UN|1|Unknown
0019|Harmony R1.0|52|UN|1|Unknown
0019|Harmony R1.0|54|UN|1|Unknown
0019|Harmony R1.0|55|UN|1|Unknown
0019|Harmony R1.0|56|US|1|Unknown
0019|Harmony R1.0|57|UN|1|Unknown
0019|Harmony R1.0|58|UN|1|Unknown
0019|Harmony R1.0|59|UN|1|Unknown
0019|Harmony R1.0|5a|UN|1|Unknown
0019|Harmony R1.0|5b|US|1|Unknown
0019|Harmony R1.0|5c|UN|1|Unknown
0019|Harmony R1.0|5d|UN|1|Unknown
0019|Harmony R1.0|5f|UI|1|Unknown
0019|Harmony R1.0|60|UI|1|Unknown
0019|Harmony R1.0|63|US|1|Unknown
0019|Harmony R1.0|64|UN|1|Unknown
0019|Harmony R1.0|65|UN|1|Unknown
0019|Harmony R1.0|66|DS|1|Unknown
0019|Harmony R1.0|67|IS|1|Unknown
0019|Harmony R1.0|68|IS|1|Unknown
0019|Harmony R1.0|69|IS|1|Unknown
0019|Harmony R1.0|6a|IS|1|Unknown
0019|Harmony R1.0|6b|LO|1|Unknown
0019|Harmony R1.0|70|LO|1|Unknown
0019|Harmony R1.0|71|LO|1|Unknown
0019|Harmony R1.0|72|IS|1|Unknown
0019|Harmony R1.0|73|IS|1|Unknown
0019|Harmony R1.0|74|US|1|Unknown
0019|Harmony R1.0|75|IS|1|Unknown
0019|Harmony R1.0|78|IS|1|Unknown
0019|Harmony R1.0|79|IS|1|Unknown
0019|Harmony R1.0|7a|IS|1|Unknown
0019|Harmony R1.0|7b|IS|1|Unknown
0019|Harmony R1.0|7c|US|1|Unknown
0019|Harmony R1.0|7d|US|1|Unknown
0019|Harmony R1.0|7e|US|1|Unknown
0019|Harmony R1.0|7f|US|1|Unknown
0019|Harmony R1.0|80|US|1|Unknown
0019|Harmony R1.0|81|US|1|Unknown
0019|Harmony R1.0|82|US|1|Unknown
0019|Harmony R1.0|83|US|1|Unknown
0019|Harmony R1.0 C2|00|LO|1|Unknown
0019|Harmony R1.0 C2|01|UN|1|Unknown
0019|Harmony R1.0 C2|02|UN|1|Unknown
0019|Harmony R1.0 C2|03|UN|1|Unknown
0019|Harmony R1.0 C2|04|UN|1|Unknown
0019|Harmony R1.0 C2|05|UN|1|Unknown
0019|Harmony R1.0 C2|06|LO|1|Unknown
0019|Harmony R1.0 C2|07|UN|1|Unknown
0019|Harmony R1.0 C2|08|UN|1|Unknown
0019|Harmony R1.0 C2|09|UN|1|Unknown
0019|Harmony R1.0 C2|0a|UN|1|Unknown
0019|Harmony R1.0 C2|6a|LO|1|Unknown
0019|Harmony R1.0 C2|6c|US|1|Unknown
0019|Harmony R1.0 C2|6d|US|1|Unknown
0019|Harmony R1.0 C2|6e|UN|1|Unknown
0019|Harmony R1.0 C2|74|UN|1|Unknown
0019|Harmony R1.0 C2|76|UN|1|Unknown
0019|Harmony R1.0 C2|78|US|1|Unknown
0019|Harmony R1.0 C2|79|US|1|Unknown
0019|Harmony R1.0 C2|7a|US|1|Unknown
0019|Harmony R1.0 C2|80|UN|1|Unknown
0019|Harmony R1.0 C2|81|UN|1|Unknown
0019|Harmony R1.0 C2|82|UN|1|Unknown
0019|Harmony R1.0 C2|83|UN|1|Unknown
0019|Harmony R1.0 C2|84|UN|1|Unknown
0019|Harmony R1.0 C2|91|UN|1|Unknown
0019|Harmony R1.0 C3|00|LO|1|Unknown
0019|Harmony R1.0 C3|03|LO|1|Unknown
0019|Harmony R1.0 C3|07|LO|1|Unknown
0019|Harmony R1.0 C3|0b|LO|1|Unknown
0019|Harmony R1.0 C3|50|UN|1|Unknown
0019|Harmony R1.0 C3|51|UN|1|Unknown
0019|Harmony R1.0 C3|52|LO|1|Unknown
0019|Harmony R1.0 C3|53|UN|1|Unknown
0019|Harmony R1.0 C3|5a|US|1|Unknown
0019|Harmony R1.0 C3|5b|LO|1|Unknown
0019|Harmony R1.0 C3|5c|US|1|Unknown
0019|Harmony R1.0 C3|5f|US|1|Unknown
0019|Harmony R1.0 C3|78|LO|1|Unknown
0019|Harmony R1.0 C3|79|PN|1|Unknown
0019|Harmony R1.0 C3|7a|PN|1|Unknown
0019|Harmony R1.0 C3|7b|LO|1|Unknown
0019|Harmony R1.0 C3|7c|UN|1|Unknown
0019|Harmony R1.0 C3|7d|CS|1|Unknown
0019|Harmony R1.0 C3|7e|LO|1|Unknown
0019|Harmony R1.0 C3|7f|UN|1|Unknown
0019|Harmony R1.0 C3|80|IS|1|Unknown
0019|Harmony R1.0 C3|83|IS|1|Unknown
0019|Harmony R1.0 C3|94|IS|1|Unknown
0019|Harmony R1.0 C3|95|IS|1|Unknown
0019|Harmony R1.0 C3|96|LO|1|Unknown
0019|Harmony R1.0 C3|97|UN|1|Unknown
0019|Harmony R1.0 C3|98|IS|1-n|Unknown
0019|Harmony R1.0 C3|e4|LO|1|Unknown
0019|Harmony R1.0 C3|e5|UN|1|Unknown
0019|Harmony R1.0 C3|e6|UN|1|Unknown
0019|Harmony R1.0 C3|e7|UN|1|Unknown
0019|Harmony R1.0 C3|e8|UN|1|Unknown
0019|Harmony R1.0 C3|e9|US|1|Unknown
0019|Harmony R1.0 C3|ea|UN|1|Unknown
0019|Harmony R1.0 C3|eb|US|1|Unknown
0019|Harmony R1.0 C3|ec|UN|1|Unknown
0019|Harmony R1.0 C3|ed|UN|1|Unknown
0019|Harmony R1.0 C3|ee|US|1|Unknown
0019|Harmony R1.0 C3|ef|US|1|Unknown
0019|Harmony R1.0 C3|f0|UN|1|Unknown
0019|Harmony R1.0 C3|f1|UN|1|Unknown
0019|Harmony R1.0 C3|f2|UN|1|Unknown
0019|Harmony R2.0|79|IS|1|Unknown
0019|Harmony R2.0|7c|IS|1|Unknown
0019|Harmony R2.0|7d|UN|1|Unknown
0019|Harmony R2.0|81|IS|1|Unknown
0019|Harmony R2.0|82|US|1|Unknown
0019|Harmony R2.0|83|US|1|Unknown
0019|Harmony R2.0|84|US|1|Unknown
0019|Harmony R2.0|85|UN|1|Unknown
0019|Harmony R2.0|86|IS|1|Unknown
0019|Harmony R2.0|87|UN|1|Unknown
0019|Harmony R2.0|88|IS|1|Unknown
0019|Harmony R2.0|89|US|1|Unknown
0019|Harmony R2.0|8a|US|1|Unknown
0019|Harmony R2.0|8c|IS|1|Unknown
0019|Harmony R2.0|8d|DS|1|Unknown
0019|Harmony R2.0|8f|US|1|Unknown
0019|Harmony R2.0|90|US|1|Unknown
0019|Harmony R2.0|91|US|1|Unknown
0019|Harmony R2.0|92|US|1|Unknown
0019|Harmony R2.0|93|DS|2|Unknown
0019|Harmony R2.0|94|LO|1|Unknown
0019|Harmony R2.0|95|LO|1-n|Unknown
0019|Harmony R2.0|96|DS|1|Unknown
0019|Harmony R2.0|97|IS|2|Unknown
0019|Harmony R2.0|99|LO|1|Unknown
0029|Silhouette V1.0|31|UN|1|Unknown
0029|Silhouette V1.0|46|UN|1|Unknown
0029|Silhouette V1.0|47|UN|1|Unknown
0029|Silhouette V1.0|73|UN|1|Unknown
0029|Silhouette V1.0|74|UN|1|Unknown
0029|Silhouette V1.0|77|UN|1|Unknown
0029|Silhouette V1.0|78|UN|1|Unknown
0029|Silhouette V1.0|88|UN|1|Unknown
0029|Silhouette V1.0|89|UN|1|Unknown
0029|Silhouette V1.0|90|UN|1|Unknown
0029|Silhouette V1.0|91|UN|1|Unknown
0011|Hologic|00|OB|1|Hx Questionnaire
0011|HOLOGIC|00|OB|1|Hx Questionnaire
0013|Hologic|00|LO|1|IVA Results Flag
0013|HOLOGIC|00|LO|1|IVA Results Flag
0019|Hologic|00|UT|1|Report Data
0019|HOLOGIC|00|UT|1|Report Data
0019|LODOX_STATSCAN|01|IS|1-n|Unknown
0019|LODOX_STATSCAN|02|IS|1|Unknown
0019|LODOX_STATSCAN|03|DS|1|Unknown
0019|LODOX_STATSCAN|04|DS|1|Unknown
0019|LODOX_STATSCAN|05|DS|1|Unknown
0019|LODOX_STATSCAN|06|DS|1|Unknown
0019|LODOX_STATSCAN|07|DS|1|Unknown
0019|LODOX_STATSCAN|08|DS|1|Unknown
0021|SCHICK TECHNOLOGIES - Change List Creator ID|01|UI|1|Unknown
0021|SCHICK TECHNOLOGIES - Change List Creator ID|02|SQ|1|Unknown
0021|SCHICK TECHNOLOGIES - Note List Creator ID|01|UI|1|Unknown
0021|SCHICK TECHNOLOGIES - Note List Creator ID|02|SQ|1|Unknown
0021|SCHICK TECHNOLOGIES - Change Item Creator ID|01|UI|1|Unknown
0021|SCHICK TECHNOLOGIES - Change Item Creator ID|02|US|1|Unknown
0021|SCHICK TECHNOLOGIES - Change Item Creator ID|03|DT|1|Unknown
0021|SCHICK TECHNOLOGIES - Change Item Creator ID|04|PN|1|Unknown
0021|SCHICK TECHNOLOGIES - Change Item Creator ID|05|OB|1|Unknown
0021|Hologic|01|LT|1|Image Analysis Data in XML
0021|HOLOGIC|01|LT|1|Image Analysis Data in XML
0023|Hologic|00|LO|1|Encoding Scheme Version
0023|HOLOGIC|00|LO|1|Encoding Scheme Version
0023|Hologic|01|LO|1|P File Name
0023|HOLOGIC|01|LO|1|P File Name
0023|Hologic|02|OB|1|P File Data
0023|HOLOGIC|02|OB|1|P File Data
0023|Hologic|03|UL|1|P File Length
0023|HOLOGIC|03|UL|1|P File Length
0023|Hologic|04|OB|1|R File Data
0023|HOLOGIC|04|OB|1|R File Data
0023|Hologic|05|UL|1|R File Length
0023|HOLOGIC|05|UL|1|R File Length
0029|Hologic|00|OB|1|Graph Bitmap Data
0029|HOLOGIC|00|OB|1|Graph Bitmap Data
0029|Hologic|01|UL|1|Graph Bitmap Size
0029|HOLOGIC|01|UL|1|Graph Bitmap Size
0029|SCHICK TECHNOLOGIES - Image Security Creator ID|01|UL|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|20|LT|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|21|ST|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|22|ST|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|23|ST|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|24|LO|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|25|LO|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|26|LO|1|Unknown
0029|2.16.840.1.114059.1.1.6.1.50.1|27|LO|1|Unknown
0073|STENTOR|01|ST|1|Unknown
0073|STENTOR|02|ST|1|Unknown
0073|STENTOR|03|ST|1|Unknown
0073|STENTOR|04|ST|1|Unknown
0073|STENTOR|06|LO|1|Unknown
0119|MRSC|1204|IS|1|NumberPasses
0019|FDMS 1.0|30|LO|1|Menu Character String
0021|FDMS 1.0|70|IS|1|Film Number within the Series
0021|FDMS 1.0|90|CS|1|LUT Number
0009|FDMS 1.0|f1|LO|1|Processing Information Flag
0019|MMCPrivate|03|SH|1|Is Snap Shot Series
0029|FDMS 1.0|25|CS|1|Image Rotation/Reversal Information
0032|FDMS 1.0|32|PN|1|Requesting Physician
0032|FDMS 1.0|33|LO|1|Requesting Service
2011|FDMS 1.0|00|CS|1|Trim Density
2011|FDMS 1.0|01|IS|1|Trim Width
2011|FDMS 1.0|02|CS|1|Image Mag./Reduc. Range
2011|FDMS 1.0|10|CS|1|Image Display Format
2011|FDMS 1.0|20|OW|1|Interpolation A-VRS System Format
50f1|FDMS 1.0|10|CS|1|Film Output Format
0019|Canon Inc.|10|UN|1|Unknown
0019|Canon Inc.|13|UN|1|Unknown
0019|Canon Inc.|15|DS|2|Unknown
0019|Canon Inc.|16|UN|1|Unknown
0019|Canon Inc.|17|DS|1|Unknown
0019|Canon Inc.|18|UN|1|Unknown
0019|Canon Inc.|19|UN|1|Unknown
0019|Canon Inc.|1a|UN|1|Unknown
0019|Canon Inc.|1b|LO|1|Unknown
0019|Canon Inc.|1c|IS|1|Unknown
0019|Canon Inc.|1e|IS|1|Unknown
0019|Canon Inc.|1f|UN|1|Unknown
0019|Canon Inc.|21|IS|1|Unknown
50f1|FDMS 1.0|0a|LO|1|FNC Parameters
0009|SECTRA_Ident_01|01|SH|1|Request number
0009|SECTRA_Ident_01|02|SH|1|Examination number
0009|SECTRA_Ident_01|04|LO|1|Series Identifier
0009|SECTRA_Ident_01|05|LO|1|Series Order
0009|SECTRA_Ident_01|06|LO|1|File Name
0009|SECTRA_Ident_01|07|LO|1|Image Data ID
0029|SECTRA_ImageInfo_01|01|OB|1|Image info
0029|SECTRA_ImageInfo_01|02|CS|1|Marking
0029|SECTRA_ImageInfo_01|03|LO|1|No decompression
0029|SECTRA_ImageInfo_01|04|OB|1|Image info new
6001|SECTRA_OverlayInfo_01|01|LO|1|Sectra Overlay
0009|BioPri|00|LO|1|Unknown
0009|BioPri|01|UN|1|Unknown
0009|BioPri|02|UN|1|Unknown
0009|BioPri|03|LO|1-n|Unknown
0009|BioPri|04|LO|1|Unknown
0009|BioPri|05|LO|1|Unknown
0009|BioPri|07|LO|1|Unknown
0009|BioPri|08|LO|1|Unknown
0009|BioPri|09|LO|1|Unknown
0009|BioPri|10|UN|1|Unknown
0029|Silhouette VRS 3.0|13|UN|1|Unknown
0029|Silhouette VRS 3.0|14|UN|1|Unknown
0029|Silhouette VRS 3.0|17|UN|1|Unknown
0029|Silhouette VRS 3.0|18|UN|1|Unknown
0029|Silhouette VRS 3.0|19|UN|1|Unknown
0029|Silhouette VRS 3.0|1a|UN|1|Unknown
0029|Silhouette VRS 3.0|1b|UN|1|Unknown
0029|Silhouette VRS 3.0|1c|UN|1|Unknown
0029|Silhouette VRS 3.0|1d|UN|1|Unknown
0019|ADAC_IMG|21|US|1|Number of ADAC Headers
0019|ADAC_IMG|41|IS|1-n|ADAC Header/Image Size
0019|ADAC_IMG|61|OB|1|ADAC Pegasys Headers
0029|Silhouette VRS 3.0|1e|UN|1|Unknown
0029|Silhouette VRS 3.0|27|US|1|Unknown
0029|Silhouette VRS 3.0|28|UN|1|Unknown
0029|Silhouette VRS 3.0|30|UN|1|Unknown
0029|Silhouette VRS 3.0|32|UN|1|Unknown
0029|Silhouette VRS 3.0|34|UN|1|Unknown
0029|Silhouette VRS 3.0|35|CS|1|Unknown
0029|Silhouette VRS 3.0|36|US|1|Unknown
0011|Hipaa Private Creator|01|LT|1|Encrypted Instance Creator ID
0011|Hipaa Private Creator|02|LT|1|Encrypted SOP Instance UID
0011|Hipaa Private Creator|03|LT|1|Encrypted Accession Number
0011|Hipaa Private Creator|04|LT|1|Encrypted Institution Name
0011|Hipaa Private Creator|05|LT|1|Encrypted Institution Address
0011|Hipaa Private Creator|06|LT|1|Encrypted Referring Physician's Name
0011|Hipaa Private Creator|07|LT|1|Encrypted Referring Physician's Address
0011|Hipaa Private Creator|08|LT|1|Encrypted Station Name
0011|Hipaa Private Creator|09|LT|1|Encrypted Study Description
0011|Hipaa Private Creator|10|LT|1|Encrypted Series Description
0011|Hipaa Private Creator|11|LT|1|Encrypted Institutional Department Name
0011|Hipaa Private Creator|12|LT|1|Encrypted Physicians of Record
0011|Hipaa Private Creator|13|LT|1|Encrypted Performing Physician's Name
0011|Hipaa Private Creator|14|LT|1|Encrypted Name of Physicians Reading Study
0011|Hipaa Private Creator|15|LT|1|Encrypted Operator's Name
0011|Hipaa Private Creator|16|LT|1|Encrypted Admitting Diagnoses Description
0011|Hipaa Private Creator|17|LT|1|Encrypted Referenced SOP Instance UID
0011|Hipaa Private Creator|18|LT|1|Encrypted Derivation Description
0011|Hipaa Private Creator|19|LT|1|Encrypted Patient's Name
0011|Hipaa Private Creator|20|LT|1|Encrypted Patient's ID
0011|Hipaa Private Creator|21|LT|1|Encrypted Patient's Birth Date
0011|Hipaa Private Creator|22|LT|1|Encrypted Patient's Birth Time
0011|Hipaa Private Creator|23|LT|1|Encrypted Patient's Sex
0011|Hipaa Private Creator|24|LT|1|Encrypted Other Patient IDs
0011|Hipaa Private Creator|25|LT|1|Encrypted Other Patient Names
0011|Hipaa Private Creator|26|LT|1|Encrypted Patient's Age
0011|Hipaa Private Creator|27|LT|1|Encrypted Patient's Size
0011|Hipaa Private Creator|28|LT|1|Encrypted Patient's Weight
0011|Hipaa Private Creator|29|LT|1|Encrypted Medical Record Locator
0011|Hipaa Private Creator|30|LT|1|Encrypted Ethnic Group
0011|Hipaa Private Creator|31|LT|1|Encrypted Occupation
0011|Hipaa Private Creator|32|LT|1|Encrypted Additional Patient's History
0011|Hipaa Private Creator|33|LT|1|Encrypted Patient Comments
0011|Hipaa Private Creator|34|LT|1|Encrypted Device Serial Number
0011|Hipaa Private Creator|35|LT|1|Encrypted Protocol Name
0011|Hipaa Private Creator|36|LT|1|Encrypted Study Instance UID
0011|Hipaa Private Creator|37|LT|1|Encrypted Series Instance UID
0011|Hipaa Private Creator|38|LT|1|Encrypted Study ID
0011|Hipaa Private Creator|39|LT|1|Encrypted Frame of Reference UID
0119|MRSC|1206|IS|1-n|NumProcesses
0011|Hipaa Private Creator|40|LT|1|Encrypted Synchronization Frame of Reference UID
0011|Hipaa Private Creator|41|LT|1|Encrypted Image Comments
0011|Hipaa Private Creator|42|LT|1|Encrypted UID
0019|LORAD Selenia|06|LO|1|Paddle ID
0019|LORAD Selenia|07|SH|1|Paddle Position
0019|LORAD Selenia|08|LO|1|Collimation Size
0019|LORAD Selenia|16|DS|1|Paddle Angle
0019|LORAD Selenia|26|LO|1|Paddle ID Description
0019|LORAD Selenia|27|SH|1|Paddle Position Description
0019|LORAD Selenia|28|LO|1|Collimation Size Description
0019|LORAD Selenia|29|LO|1|AEC User Density Scale Factor Description
0019|LORAD Selenia|30|US|1|AEC User Density Scale Factor
0019|LORAD Selenia|31|US|1|AEC System Density Scale Factor
0019|LORAD Selenia|32|US|1|AEC Calculated mAs
0019|LORAD Selenia|33|US|1|AEC Auto Pixel 1
0019|LORAD Selenia|34|US|1|AEC Auto Pixel 2
0019|LORAD Selenia|35|US|1|AEC Sensor
0019|LORAD Selenia|37|LO|1|NPT Mode
0019|LORAD Selenia|40|DS|1|Skin Edge
0019|LORAD Selenia|41|DS|1|Exposure Index
0019|LORAD Selenia|50|DS|1|Display Minimum OD
0019|LORAD Selenia|51|DS|1|Dispaly Maximum OD
0019|LORAD Selenia|52|IS|1|Display Minimum Nits
0019|LORAD Selenia|53|IS|1|Display Maximum Nits
0019|LORAD Selenia|60|LT|1|Geometry Calibration
0019|LORAD Selenia|70|LO|1|Frame of Reference ID
0019|LORAD Selenia|71|CS|1|Paired Position
0019|LORAD Selenia|80|SH|1|Detector Image Offset
0019|LORAD Selenia|90|DS|1|Conventional Tomo Angle
0019|HOLOGIC, Inc.|01|IS|1|Unknown
0019|HOLOGIC, Inc.|02|IS|1|Unknown
0019|HOLOGIC, Inc.|03|IS|1|Unknown
0019|HOLOGIC, Inc.|04|IS|1|Unknown
0019|HOLOGIC, Inc.|06|LO|1|Paddle ID
0019|HOLOGIC, Inc.|07|SH|1|Paddle Position
0019|HOLOGIC, Inc.|08|LO|1|Collimation Size
0019|HOLOGIC, Inc.|16|DS|1|Paddle Angle
0019|HOLOGIC, Inc.|25|SH|1|Unknown
0019|HOLOGIC, Inc.|26|LO|1|Paddle ID Description
0019|HOLOGIC, Inc.|27|SH|1|Paddle Position Description
0019|HOLOGIC, Inc.|28|LO|1|Collimation Size Description
0019|HOLOGIC, Inc.|29|LO|1|AEC User Density Scale Factor Description
0019|HOLOGIC, Inc.|30|US|1|AEC User Density Scale Factor
0019|HOLOGIC, Inc.|31|US|1|AEC System Density Scale Factor
0019|HOLOGIC, Inc.|32|US|1|AEC Calculated mAs
0019|HOLOGIC, Inc.|33|US|1|AEC Auto Pixel 1
0019|HOLOGIC, Inc.|34|US|1|AEC Auto Pixel 2
0019|HOLOGIC, Inc.|35|US|1|AEC Sensor
0019|HOLOGIC, Inc.|37|LO|1|NPT Mode
0019|HOLOGIC, Inc.|40|DS|1|Skin Edge
0019|HOLOGIC, Inc.|41|DS|1|Exposure Index
0019|HOLOGIC, Inc.|42|IS|1|Exposure Index Target
0019|HOLOGIC, Inc.|43|DS|1|Short Index Ratio
0019|HOLOGIC, Inc.|44|DS|1|Scout kVp
0019|HOLOGIC, Inc.|45|IS|1|Scout mA
0019|HOLOGIC, Inc.|46|IS|1|Scout mAs
0019|HOLOGIC, Inc.|50|DS|1|Display Minimum OD
0019|HOLOGIC, Inc.|51|DS|1|Dispaly Maximum OD
0019|HOLOGIC, Inc.|52|IS|1|Display Minimum Nits
0019|HOLOGIC, Inc.|53|IS|1|Display Maximum Nits
0019|HOLOGIC, Inc.|60|LT|1|Geometry Calibration
0019|HOLOGIC, Inc.|61|OB|1|3D IP Parameters
0019|HOLOGIC, Inc.|62|LT|1|2D IP Parameters
0019|HOLOGIC, Inc.|70|LO|1|Frame of Reference ID
0019|HOLOGIC, Inc.|71|CS|1|Paired Position
0019|HOLOGIC, Inc.|80|SH|1|Detector Image Offset
0019|HOLOGIC, Inc.|85|SH|1|Image Source
0019|HOLOGIC, Inc.|87|LO|1|Marker Text
0019|HOLOGIC, Inc.|88|LO|1|Marker Tech Initials
0019|HOLOGIC, Inc.|89|DS|2|Marker Location
0019|HOLOGIC, Inc.|8a|SQ|2|Marker Sequence
0019|HOLOGIC, Inc.|90|DS|1|Conventional Tomo Angle
0019|HOLOGIC, Inc.|97|SH|1|Markers Burned Into Image
0019|HOLOGIC, Inc.|98|LO|1|Grid Line Correction
7e01|HOLOGIC, Inc.|01|LO|1|Codec Version
7e01|HOLOGIC, Inc.|02|SH|1|Codec Content Type
7e01|HOLOGIC, Inc.|10|SQ|1|High Resolution Data Sequence
7e01|HOLOGIC, Inc.|11|SQ|1|Low Resolution Data Sequence
7e01|HOLOGIC, Inc.|12|OB|1|Codec Content
7f01|HOLOGIC, Inc.|01|LO|1|Codec Version
7f01|HOLOGIC, Inc.|02|SH|1|Codec Content Type
7f01|HOLOGIC, Inc.|10|SQ|1|High Resolution Data Sequence
7f01|HOLOGIC, Inc.|11|SQ|1|Low Resolution Data Sequence
7f01|HOLOGIC, Inc.|12|OB|1|Codec Content
0029|1.2.840.113663.1|00|US|1|Unknown
0029|1.2.840.113663.1|01|US|1|Unknown
0009|MMCPrivate|50|CS|1|CMS Patient Position
0009|MMCPrivate|51|LO|1|CMI Contrast Bolus Agent
0009|MMCPrivate|52|LO|1|CMS institution Name
0009|MMCPrivate|53|LO|1|CMS Institutional Department Name
0009|MMCPrivate|54|LO|1|CMS Series Description
0009|MMCPrivate|55|LO|1|CMS Operators Name
0009|MMCPrivate|56|LO|1|CMS Performing Physicians Name
0009|MMCPrivate|57|ST|1|CMS Institution Address
0009|MMCPrivate|58|LO|1|CMI Image Comments
0009|MMCPrivate|59|LO|1|CMI Instance Creation DateTime
0009|MMCPrivate|5a|LO|1|MPPS Step Status
0009|MMCPrivate|5b|IS|1|Filmed Count
0009|MMCPrivate|5c|LO|1|Is Allow Cascade Save
0009|MMCPrivate|5d|LO|1|Is Allow Cascade Protect
0009|MMCPrivate|5e|LO|1|Is Deleted
0011|MMCPrivate|03|IS|1|Filmed Count
0011|MMCPrivate|04|OB|1|Application Data
0011|MMCPrivate|05|LO|1|Is Allow Cascade Save
0011|MMCPrivate|06|LO|1|Is Allow Cascade Protect
0011|MMCPrivate|07|LO|1|Is Deleted
0009|MMCPrivate|02|LO|1|Scheduled Study DateTime
0009|MMCPrivate|03|OB|1|Study App Data
0009|MMCPrivate|48|LO|1|Protocol Name
0009|MMCPrivate|4e|LO|1|CMS Body Part Examined
0009|MMCPrivate|4f|LO|1|Is Protected
0011|MMCPrivate|01|LO|1|Is Rapid Registration
0011|MMCPrivate|02|LO|1|Is Protected
0019|MMCPrivate|01|LO|1|Proc Type
0019|MMCPrivate|02|LO|1|Plane
0119|MRSC|1208|IS|1-n|GroupExecuteOrder
0019|MMCPrivate|12|IS|1|Image Increment
0019|MMCPrivate|13|LO|1|MPPS Step Status
0019|MMCPrivate|14|IS|1|Storage Committed Count
0019|MMCPrivate|15|IS|1|Archived Count
0019|MMCPrivate|16|IS|1|Transferred Count
0019|MMCPrivate|17|LO|1|Is Allow Cascade Save
0019|MMCPrivate|18|LO|1|Is Allow Cascade Protect
0019|MMCPrivate|19|LO|1|Is Deleted
0019|MMCPrivate|1a|UI|1|Characterized Image Instance UID
0019|MMCPrivate|1b|IS|1|Characterized Image Count
0019|MMCPrivate|1c|LO|1|Internal Window Width
0019|MMCPrivate|1d|LO|1|Internal Window Level
0019|MMCPrivate|1e|LO|1|Unknown
0019|MMCPrivate|07|LO|1|Image Contrast Bolus Agent
0019|MMCPrivate|08|DS|1|Image Slice Thickness
0019|MMCPrivate|0a|LO|1|Image Echo Time
0019|MMCPrivate|0b|DS|1|Image Repetition Time
0019|MMCPrivate|0c|LO|1|Sequence Type
0019|MMCPrivate|0d|LO|1|Task UID
0019|MMCPrivate|0e|OB|1|Series App Data
0019|MMCPrivate|0f|IS|1|Multi Slice Number
0019|MMCPrivate|10|LO|1|Image Scan Time
0019|MMCPrivate|11|LO|1|Is Protected
0029|MMCPrivate|01|IS|1|Slice Number
0029|MMCPrivate|02|IS|1|Phase Number
0029|MMCPrivate|03|LO|1|Proc Type
0029|MMCPrivate|04|LO|1|Stopwatch Time
0029|MMCPrivate|05|LO|1|Plane
0029|MMCPrivate|06|LO|1|Scan Time
0029|MMCPrivate|08|LO|1|Dual Slice Flag
0029|MMCPrivate|09|LO|1|SSP Ratio
0029|MMCPrivate|0a|LO|1|Gating Signal Source
0029|MMCPrivate|0b|LO|1|Rephase
0029|MMCPrivate|0c|LO|1|Half Echo
0029|MMCPrivate|0d|LO|1|Rect FOV Ratio
0029|MMCPrivate|0e|LO|1|Half Scan
0029|MMCPrivate|0f|LO|1|Num Shots
0029|MMCPrivate|10|LO|1|Contrast Agent
0029|MMCPrivate|12|LO|1|Num Echo Shift
0029|MMCPrivate|13|LO|1|Fat Sat
0029|MMCPrivate|14|LO|1|MTC
0029|MMCPrivate|15|LO|1|Num Pre Sat
0029|MMCPrivate|16|LO|1|Target Velocity
0029|MMCPrivate|17|LO|1|VENC Axis
0029|MMCPrivate|18|LO|1|Num VENC Direction
0029|MMCPrivate|1c|LO|1|Is Scalable Window Level
0029|MMCPrivate|1d|LO|1|Three D Setting Line Angle
0029|MMCPrivate|1e|LO|1|MPG Total Axis
0029|MMCPrivate|1f|LO|1|MPG Axis Number
0029|MMCPrivate|20|IS|1|Multi Echo Number
0029|MMCPrivate|21|DS|1|Navi Average Gate Width
0029|MMCPrivate|22|ST|1|Shim Compensate Value
0029|MMCPrivate|23|LO|1|GC Offset
0029|MMCPrivate|24|DS|1|Navi Max Gate Width
0029|MMCPrivate|25|DS|1|Navi Min Gate Width
0029|MMCPrivate|26|DS|1|Navi Max Gate Position
0029|MMCPrivate|27|DS|1|Navi Min Gate Position
0029|MMCPrivate|28|DS|1|Time Duration
0029|MMCPrivate|2a|DS|1|Navi Initial Gate Width
0119|MRSC|120a|IS|1|NumberTransforms
0029|MMCPrivate|2c|DS|1|Navi Initial Gate Position
0029|MMCPrivate|2e|DS|1|Navi Average Gate Position
0029|MMCPrivate|2f|OB|1|Image App Data
0029|MMCPrivate|30|FD|1|Diffusion BValue
0029|MMCPrivate|31|SQ|1|Shared Functional Groups Sequence
0029|MMCPrivate|32|SQ|1|Per Frame Functional Groups Sequence
0029|MMCPrivate|33|DS|1|Lossy Image Compression Ratio
0029|MMCPrivate|34|UI|1|Instance Creator UID
0029|MMCPrivate|35|UI|1|Related General SOPClass UID
0029|MMCPrivate|36|UI|1|Original Specialized SOPClass UID
0029|MMCPrivate|37|SH|1|Timezone Offset From UTC
0029|MMCPrivate|38|CS|1|SOPInstance Status
0029|MMCPrivate|39|DT|1|SOPAuthorization Dateand Time
0029|MMCPrivate|3a|LT|1|SOPAuthorization Comment
0029|MMCPrivate|3b|LO|1|Authorization Equipment Certification Number
0029|MMCPrivate|3c|UL|1|Concatenation Frame Offset Number
0029|MMCPrivate|3d|US|1|Representative Frame Number
0029|MMCPrivate|3e|UI|1|Concatenation UID
0029|MMCPrivate|3f|US|1|In Concatenation Number
0029|MMCPrivate|40|CS|1|Cardiac Synchronization Technique
0029|MMCPrivate|41|CS|1|Cardiac Signal Source
0029|MMCPrivate|42|FD|1|Cardiac RRInterval Specified
0029|MMCPrivate|43|CS|1|Cardiac Beat Rejection Technique
0029|MMCPrivate|44|IS|1|Low RR Value
0029|MMCPrivate|45|IS|1|High RR Value
0029|MMCPrivate|46|IS|1|Intervals Acquired
0029|MMCPrivate|47|IS|1|Intervals Rejected
0029|MMCPrivate|49|CS|1|Respiratory Signal Source
0029|MMCPrivate|4a|CS|1|Bulk Motion Compensation Technique
0029|MMCPrivate|4b|CS|1|Bulk Motion Signal Source
0029|MMCPrivate|4c|CS|1|Pixel Presentation
0029|MMCPrivate|4d|CS|1|Volumetric Properties
0029|MMCPrivate|4e|CS|1|Volume Based Calculation Technique
0029|MMCPrivate|4f|ST|1|Acquisition Context Description
0029|MMCPrivate|50|SQ|1|Unknown
0029|MMCPrivate|51|LO|1|LUTDescriptor
0029|MMCPrivate|52|LO|1|LUTExplanation
0029|MMCPrivate|53|LO|1|LUTData
0029|MMCPrivate|54|CS|1|Presentation LUT Shape
0029|MMCPrivate|55|SQ|1|Frame Anatomy Sequence
0029|MMCPrivate|56|CS|1|Frame Laterality
0029|MMCPrivate|57|SQ|1|Anatomic Region Sequence
0029|MMCPrivate|58|SH|1|Anatomic Region Code Value
0029|MMCPrivate|59|SH|1|Anatomic Region Coding Scheme Designator
0029|MMCPrivate|5a|SH|1|Anatomic Region Coding Scheme Version
0029|MMCPrivate|5b|LO|1|Anatomic Region Code Meaning
0029|MMCPrivate|5c|SQ|1|Pixel Value Transformation Sequence
0029|MMCPrivate|5d|LO|1|Rescale Type
0029|MMCPrivate|5e|SQ|1|Cardiac Synchronization Sequence
0029|MMCPrivate|5f|FD|1|Trigger Delay Time
0029|MMCPrivate|60|SQ|1|Frame VOILUTSequence
0029|MMCPrivate|62|CS|1|Unknown
0029|MMCPrivate|63|SQ|1|MRModifier Sequence
0029|MMCPrivate|64|CS|1|Parallel Acquisition Technique
0029|MMCPrivate|65|FD|1|Parallel Reduction Factor Sec In
0119|MRSC|120b|IS|1-n|NumberProcesses
0029|MMCPrivate|67|CS|1|Flow Compensation
0029|MMCPrivate|68|CS|1|Flow Compensation Direction
0029|MMCPrivate|69|CS|1|Spatial PreSaturation
0029|MMCPrivate|6b|CS|1|Partial Fourier Direction
0029|MMCPrivate|70|SQ|1|MR Receive Coil Sequence
0029|MMCPrivate|71|LO|1|Receive Coil Manufacturer Name
0029|MMCPrivate|72|CS|1|Receive Coil Type
0029|MMCPrivate|73|CS|1|Quadrature Receive Coil
0029|MMCPrivate|74|LO|1|Multi Coil Configuration
0029|MMCPrivate|75|CS|1|Complex Image Component
0029|MMCPrivate|76|SH|1|Pulse Sequence Name
0029|MMCPrivate|77|CS|1|Echo Pulse Sequence
0029|MMCPrivate|78|CS|1|Multiple Spin Echo
0029|MMCPrivate|79|CS|1|Multi Planar Excitation
0029|MMCPrivate|7a|CS|1|Phase Contrast
0029|MMCPrivate|7b|CS|1|Time of Flight Contrast
0029|MMCPrivate|7c|CS|1|Steady State Pulse Sequence
0029|MMCPrivate|7d|CS|1|Echo Planar Pulse Sequence
0029|MMCPrivate|7e|CS|1|Spectrally Selected Suppression
0029|MMCPrivate|7f|CS|1|Oversampling Phase
0029|MMCPrivate|80|CS|1|Segmented KSpace Traversal
0029|MMCPrivate|81|CS|1|Coverage of KSpace
0029|MMCPrivate|82|SQ|1|MR Timing and Related Parameters Sequence
0029|MMCPrivate|83|US|1|RF Echo Train Length
0029|MMCPrivate|84|US|1|Gradient Echo Train Length
0029|MMCPrivate|85|CS|1|Gradient Output Type
0029|MMCPrivate|86|FD|1|Gradient Output
0029|MMCPrivate|87|SQ|1|MRFOVGeometry Sequence
0029|MMCPrivate|89|US|1|MRAcquisition Phase Encoding Steps In Plane
0029|MMCPrivate|8a|US|1|MRAcquisitionPhase Encoding Steps Out of Plane
0029|MMCPrivate|8b|SQ|1|MR Transmit Coil Sequence
0029|MMCPrivate|8c|SH|1|Transmit Coil Name
0029|MMCPrivate|8d|LO|1|Transmit Coil Manufacturer Name
0029|MMCPrivate|8e|CS|1|Transmit Coil Type
0029|MMCPrivate|8f|SQ|1|MR Echo Sequence
0029|MMCPrivate|90|FD|1|Effective Echo Time
0029|MMCPrivate|91|SQ|1|MR Metabolite Map Sequence
0029|MMCPrivate|92|ST|1|Metabolite Map Description
0029|MMCPrivate|93|SQ|1|Metabolite Map Code Sequence
0029|MMCPrivate|94|SH|1|Metabolite Map Code Value
0029|MMCPrivate|95|SH|1|Metabolite Map Coding Scheme Designator
0029|MMCPrivate|96|SH|1|Metabolite Map Coding Scheme Version
0029|MMCPrivate|97|LO|1|Metabolite Map Code Meaning
0029|MMCPrivate|98|SQ|1|MR Imaging Modifier Sequence
0029|MMCPrivate|99|CS|1|Magnetization Transfer
0029|MMCPrivate|9a|CS|1|Blood Signal Nulling
0029|MMCPrivate|9b|CS|1|Tagging
0029|MMCPrivate|9c|FD|1|Tag Spacing First Dimension
0029|MMCPrivate|9d|FD|1|Tag Spacing Second Dimension
0029|MMCPrivate|9e|FD|1|Tag Angle First Axis
0029|MMCPrivate|9f|SS|1|Tag Angle Second Axis
0029|MMCPrivate|a0|FD|1|Tag Thickness
0029|MMCPrivate|a1|FD|1|Tagging Delay
0029|MMCPrivate|a3|DS|1|Pixel Bandwidth
0029|MMCPrivate|a4|SQ|1|MRVelocity Encoding Sequence
0119|MRSC|1211|IS|1-n|InvertImage
0029|MMCPrivate|ad|IS|1|Filmed Count
0029|MMCPrivate|ae|LO|1|Is Transferred
0029|MMCPrivate|af|LO|1|Is Archived
0029|MMCPrivate|b0|LO|1|MPPS Step Status
0029|MMCPrivate|b1|LO|1|Commitment Status
0029|MMCPrivate|b2|LO|1|Is Storage Committed
0029|MMCPrivate|b3|LO|1|Is Dicom
0029|MMCPrivate|b4|LO|1|Is Allow Cascade Save
0029|MMCPrivate|b5|LO|1|Is Allow Cascade Protect
0029|MMCPrivate|b6|LO|1|Is Deleted
0029|MMCPrivate|b7|OB|1|Application Data
0029|MMCPrivate|b8|LO|1|Is Allow Cascade Save
0029|MMCPrivate|b9|LO|1|Is Allow Cascade Protect
0029|MMCPrivate|ba|LO|1|Is Deleted
0029|MMCPrivate|bb|IS|1|VOI 1
0029|MMCPrivate|bc|IS|1|VOI 2
0029|MMCPrivate|c0|FD|1|Selective IR Column
0019|MeVis BreastCare|01|LO|1|Annotation Version
0071|MeVis BreastCare|01|LO|1|XML Formatted Text Value
0065|Viewing Protocol|93|CS|1|Unknown
1455|Mortara_Inc|00|OW|1|ELI Interpretation Vector
1455|Mortara_Inc|01|UN|1|Custom ID
1455|Mortara_Inc|02|UT|1|Race
1455|Mortara_Inc|03|UT|1|Social Security Number
1455|Mortara_Inc|04|UT|1|Attending Physician
1455|Mortara_Inc|05|UT|1|Procedural Diagnosis
1455|Mortara_Inc|06|UT|1|Note 1
1455|Mortara_Inc|07|UT|1|Note 2
1455|Mortara_Inc|08|LO|1|Order Request Number
1455|Mortara_Inc|10|LO|1|Manufacturer Name
0029|SEGAMI_HEADER|31|CS|1|Unknown
0029|SEGAMI_HEADER|32|OW|1|Unknown
0031|SEGAMI MIML|98|OW|1|Unknown
0033|SEGAMI__PAGE|97|IS|1|Unknown
0033|SEGAMI__PAGE|98|OW|1|Unknown
0035|SEGAMI__MEMO|97|SH|1|Unknown
0035|SEGAMI__MEMO|98|LT|1|Unknown
5473|MedIns HP Extensions|03|LO|1|Unknown
0029|MEDIFACE|01|UL|1|Unknown
0029|MEDIFACE|10|DS|1|Unknown
0029|MEDIFACE|11|DS|1|Unknown
0029|MMCPrivate|a6|FD|1|Velocity Encoding Minimum Value
0029|MMCPrivate|a7|FD|1|Velocity Encoding Maximum Value
0029|MMCPrivate|a8|SQ|1|MR Image Frame Type Sequence
0029|MMCPrivate|a9|CS|1|Frame Type
0029|MMCPrivate|aa|CS|1|Pixel Presentation
0029|MMCPrivate|ac|CS|1|Volume Based Calculation Technique
0029|MMCPrivate|bd|DS|1|Mixing Time
0029|MMCPrivate|be|FD|1|Selective IR Position
0029|MMCPrivate|bf|FD|1|Selective IR Row
0029|MMCPrivate|c1|FD|1|Selective IR Orientation
0029|MMCPrivate|c2|DS|1|Selective IR Thickness
0029|MMCPrivate|c3|CS|1|Rephase Order Slice
0029|MMCPrivate|c4|CS|1|Rephase Order Phase
0029|MMCPrivate|c5|CS|1|Rephase Order Freq
0029|MMCPrivate|d0|LO|1|Unknown
0029|MMCPrivate|d3|LO|1|Unknown
0029|MMCPrivate|d5|UI|1|Unknown
0029|MMCPrivate|d6|LO|1|Unknown
0029|MMCPrivate|d7|OB|1|Unknown
0029|MEDIFACE|20|DS|1|Unknown
0029|MEDIFACE|21|UL|1|Unknown
0029|MEDIFACE|22|DS|2|Unknown
0029|MEDIFACE|30|LT|1|Unknown
8003|Image (ID, Version, Size, Dump, GUID)|00|LO|1|ID
8003|Image (ID, Version, Size, Dump, GUID)|10|LO|1|Version
8003|Image (ID, Version, Size, Dump, GUID)|20|UL|1|Size
8003|Image (ID, Version, Size, Dump, GUID)|30|OB|1|Dump
8003|Image (ID, Version, Size, Dump, GUID)|40|LO|1|GUID
8101|ObjectModel (ID, Version, Place, PlaceDescription)|00|LO|1|ID
8101|ObjectModel (ID, Version, Place, PlaceDescription)|10|LO|1|Version
0015|INFINITT_FMX|10|LO|1|Unknown
0015|INFINITT_FMX|11|LO|1|Unknown
0009|BrainLAB_Conversion|01|LO|1|Export Platform Name
0009|BrainLAB_Conversion|02|OB|1|Export Platform Data
3273|BrainLAB_PatientSetup|00|DS|3|Isocenter Position
3273|BrainLAB_PatientSetup|01|CS|1|Patient Position
3411|BrainLAB_BeamProfile|01|SQ|1|Beam Profile Sequence
3411|BrainLAB_BeamProfile|02|IS|1|Beam Profile Number
3411|BrainLAB_BeamProfile|03|SQ|1|Beam Parameter Sequence
3411|BrainLAB_BeamProfile|04|UT|1|Parameter Description
3411|BrainLAB_BeamProfile|05|OB|1|Parameter Data
3411|BrainLAB_BeamProfile|06|IS|1|Referenced Beam Profile Number
0011|V1|01|OB|1|User Data
0011|V1|02|DS|1|Normalization Coefficient
0011|V1|03|DS|1-n|Receiving Gain
0011|V1|04|DS|1|Mean Image Noise
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|00|UI|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|01|OB|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|02|SQ|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|06|UL|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|07|UI|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|08|SQ|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|09|UI|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|10|IS|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|13|LO|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|14|UN|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|16|LO|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|17|UN|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|18|UN|1|Unknown
1135|Voxar 2.16.124.113543.6003.1999.12.20.12.5.0|21|UL|1|Unknown
0029|Kodak Image Information|15|LO|1|Unknown
0029|Kodak Image Information|16|LO|1|Unknown
0029|Kodak Image Information|17|LO|1|Unknown
0029|Kodak Image Information|18|UT|1|Unknown
0199|NQLeft|12|FL|1|Left Nucleus Accumbens
0029|Kodak Image Information|19|IS|1|Unknown
0029|Kodak Image Information|1a|IS|1|Unknown
0037|MAROTECH Inc.|01|LO|1|Unknown
0037|MAROTECH Inc.|21|US|1|Unknown
0037|MAROTECH Inc.|22|US|1|Unknown
0037|MAROTECH Inc.|23|OB|1|Unknown
0021|BRIT Systems, Inc.|00|SQ|1|Person Information Sequence
0021|BRIT Systems, Inc.|01|LO|1|Person ID
0021|BRIT Systems, Inc.|02|PN|1|Person Name
0021|BRIT Systems, Inc.|03|LO|1|Person Role
0021|BRIT Systems, Inc.|04|SH|1|Person Home Phone
0021|BRIT Systems, Inc.|05|SH|1|Person Work Phone
0021|BRIT Systems, Inc.|06|SH|1|Person Cell Phone
0021|BRIT Systems, Inc.|07|SH|1|Person Pager Phone
0021|BRIT Systems, Inc.|08|SH|1|Person Fax Phone
0021|BRIT Systems, Inc.|09|LO|1|Person EMail
0021|BRIT Systems, Inc.|0a|ST|1|Person Address
0021|BRIT Systems, Inc.|0b|LO|1|Person Password
0021|BRIT Systems, Inc.|0c|SH|1|Person Emergency Phone
0021|BRIT Systems, Inc.|0d|LO|1|Physician ID
0021|BRIT Systems, Inc.|11|LO|1|Original Patient ID
0021|BRIT Systems, Inc.|12|UI|1|Original Study Instance UID
0021|BRIT Systems, Inc.|13|UI|1|Original Series Instance UID
0021|BRIT Systems, Inc.|14|LO|1|Master Accession Number
0021|BRIT Systems, Inc.|15|LO|1|Order Category
0021|BRIT Systems, Inc.|16|LO|1|Patient ICN
0021|BRIT Systems, Inc.|17|LO|1|Patient DFS
0021|BRIT Systems, Inc.|18|LO|1|Patient Class
0021|BRIT Systems, Inc.|19|LO|1|Patient Type
0021|BRIT Systems, Inc.|1f|LT|1|Generic String
0021|BRIT Systems, Inc.|20|LO|1|QC Study Assigned By
0021|BRIT Systems, Inc.|21|LO|1|QC Study Split By
0021|BRIT Systems, Inc.|22|LO|1|QC Study Moved By
0021|BRIT Systems, Inc.|23|LO|1|QC Study Edited By
0021|BRIT Systems, Inc.|24|LO|1|QC Series Split By
0021|BRIT Systems, Inc.|25|LO|1|QC Series Moved By
0021|BRIT Systems, Inc.|26|LO|1|QC Series Edited By
0021|BRIT Systems, Inc.|27|LO|1|QC Image Moved By
0021|BRIT Systems, Inc.|28|LO|1|QC Image Edited By
0021|BRIT Systems, Inc.|30|LO|1|QC Done Time
0021|BRIT Systems, Inc.|31|LO|1|QC Last Modification Time
0021|BRIT Systems, Inc.|32|LO|1|QC Image Accepted By
0021|BRIT Systems, Inc.|33|LO|1|QC Image Rejected By
0021|BRIT Systems, Inc.|34|DA|1|QC Done Date
0021|BRIT Systems, Inc.|50|LO|1|QC Deletion Requested
0021|BRIT Systems, Inc.|90|AE|1|Original Sender AE Title
0021|BRIT Systems, Inc.|91|LO|1|Software Title
0021|BRIT Systems, Inc.|92|SH|1|Software Version
0021|BRIT Systems, Inc.|93|LO|1|Serial Number
0021|BRIT Systems, Inc.|a0|SQ|1|Object Action Sequence
0021|BRIT Systems, Inc.|a1|ST|1|Object Action
0021|BRIT Systems, Inc.|a2|DA|1|Object Action Date
0021|BRIT Systems, Inc.|a3|TM|1|Object Action Time
0021|BRIT Systems, Inc.|a5|AE|1|Local AE Title
0021|BRIT Systems, Inc.|a6|SH|1|Local IP Address
0021|BRIT Systems, Inc.|a7|AE|1|Remote AE Title
0021|BRIT Systems, Inc.|a8|SH|1|Remote IP Address
3005|MDS NORDION OTP ANATOMY MODELLING|00|SQ|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|02|CS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|04|DS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|06|DS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|08|DS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|0a|CS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|0c|CS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|0e|CS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|10|DS|1|Unknown
3005|MDS NORDION OTP ANATOMY MODELLING|12|DS|1|Unknown
4321|Imaging Dynamics Company Ltd.|41|CS|1|Unknown
4321|Imaging Dynamics Company Ltd.|42|US|1|Unknown
4321|Imaging Dynamics Company Ltd.|64|LO|1|POD Mode
f001|Sound Technologies|00|LO|1|Patient Species
f001|Sound Technologies|01|LO|1|Patient Breed
f001|Sound Technologies|02|LO|1|Patient Category Size
f001|Sound Technologies|03|CS|1|Patient Sex Extended
f001|Sound Technologies|04|LO|1|Image View
f001|Sound Technologies|05|LO|1|Anatomy Imaged
f001|Sound Technologies|06|LT|1|Image Enhancements
f001|Sound Technologies|07|LO|1|Detector Settings
f001|Sound Technologies|08|LO|1|Application Version
f001|Sound Technologies|09|LO|1|Image Laterality Extended
f001|Sound Technologies|0a|PN|1|Client Name
f001|Sound Technologies|0b|UI|1|Reference Study Instance UID
f001|Sound Technologies|0c|UI|1|Reference Study Instance UID
f001|Sound Technologies|0d|LO|1|Exam Ref ID
f001|Sound Technologies|0e|ST|1|Physician of Record Address
f001|Sound Technologies|0f|SH|1|Physician of Record Phone Numbers
f001|Sound Technologies|10|LT|1|Reason For Study
f001|Sound Technologies|11|LO|1|Protocol
f001|Sound Technologies|12|LO|1|Capture Input Type
f001|Sound Technologies|13|LT|1|Exam Complaint
f001|Sound Technologies|14|LO|1|Exam Web Code
f001|Sound Technologies|15|LO|1|Exam Category
f001|Sound Technologies|16|SH|1|Exam Diagnosis
f001|Sound Technologies|17|PN|1|Exam Created By
f001|Sound Technologies|18|LO|1|Exam Created By Group
f001|Sound Technologies|19|DT|1|Exam Required By DateTime
f001|Sound Technologies|1a|LO|1|Capture Type
f001|Sound Technologies|1b|IS|1|Telemed Exam ID
f001|Sound Technologies|1c|LO|1|Exam Created By Guid
f001|Sound Technologies|1d|LO|1|Client Name Guid
f001|Sound Technologies|1e|LO|1|Receptor Bits Per Pixel
3711|A.L.I. Technologies, Inc.|01|LO|1|Filename
3711|A.L.I. Technologies, Inc.|02|OB|1|Data Blob of a Visit
3711|A.L.I. Technologies, Inc.|03|US|1|Revision Number
3711|A.L.I. Technologies, Inc.|04|UL|1|Unix Timestamp
3711|A.L.I. Technologies, Inc.|05|IS|1|Bag ID
3711|A.L.I. Technologies, Inc.|0c|UI|1|Original Study UID
3711|A.L.I. Technologies, Inc.|0d|US|1|Overlay Grayscale Value
3711|A.L.I. Technologies, Inc.|0e|CS|1|Anonymization Status
3711|A.L.I. Technologies, Inc.|0f|CS|1|Instance Type
3711|A.L.I. Technologies, Inc.|30|LO|1|IP Converted Frame
3711|A.L.I. Technologies, Inc.|97|OB|1|Unknown
7777|NUD_PRIVATE|02|UT|1|Interfile
7777|NUD_PRIVATE|05|IS|1|Unknown
0011|IDEXX|00|LO|1|Breed Name
0011|IDEXX|01|LO|1|Species Name
0011|IDEXX|02|PN|1|Owner
0009|WG12 Supplement 43|01|SQ|1|Event Timer Sequence
0009|WG12 Supplement 43|02|FD|1|Event Time Interval
0009|WG12 Supplement 43|03|SQ|1|Event Code Sequence
0019|WG12 Supplement 43|01|FD|1|Focus Depth(s)
0019|WG12 Supplement 43|03|SQ|1|Excluded Intervals Sequence
0019|WG12 Supplement 43|04|DT|1|Exclusion Start Datetime
0019|WG12 Supplement 43|05|FD|1|Exclusion Duration
0019|WG12 Supplement 43|06|SQ|1|US Image Description Sequence
0019|WG12 Supplement 43|07|SQ|1|Image Data Type Sequence
0019|WG12 Supplement 43|08|CS|1|Data Type
0019|WG12 Supplement 43|09|SQ|1|Transducer Scan Geometry Code Sequence
0019|WG12 Supplement 43|0b|CS|1|Aliased Data Type
0019|WG12 Supplement 43|0c|CS|1|Position Measuring Device Used
0019|WG12 Supplement 43|0d|SQ|1|Transducer Scanning Configuration Code Sequence
0019|WG12 Supplement 43|0e|SQ|1|Transducer Beam Steering Code Sequence
0019|WG12 Supplement 43|0f|SQ|1|Transducer Access Code Sequence
0021|WG12 Supplement 43|01|FD|1|Image Position (Volume)
0021|WG12 Supplement 43|02|FD|1|Image Orientation (Volume)
0021|WG12 Supplement 43|07|CS|1|Ultrasound Acquisition Geometry
0021|WG12 Supplement 43|08|FD|1|Apex Position
0021|WG12 Supplement 43|09|FD|1|Volume to Transducer Mapping Matrix
0021|WG12 Supplement 43|0a|FD|1|Volume to Table Mapping Matrix
0021|WG12 Supplement 43|0c|CS|1|Patient Frame of Reference Source
0021|WG12 Supplement 43|0d|FD|1|Temporal Position Time Offset
0021|WG12 Supplement 43|0e|SQ|1|Plane Position (Volume) Sequence
0021|WG12 Supplement 43|0f|SQ|1|Plane Orientation (Volume) Sequence
0021|WG12 Supplement 43|10|SQ|1|Temporal Position Sequence
0021|WG12 Supplement 43|11|CS|1|Dimension Organization Type
0029|WG12 Supplement 43|01|SQ|1|Data Frame Assignment Sequence
0029|WG12 Supplement 43|02|CS|1|Data Path Assignment
0029|WG12 Supplement 43|03|US|1|Bits Mapped to Color Lookup Table
0029|WG12 Supplement 43|04|SQ|1|Opacity 1 LUT Sequence
0029|WG12 Supplement 43|05|CS|1|Opacity 1 LUT Transfer Function
0029|WG12 Supplement 43|06|FD|1|Opacity Constant
0029|WG12 Supplement 43|07|US|1|Opacity Lookup Table Descriptor
0199|NQLeft|13|FL|1|Left Brain Stem
0029|WG12 Supplement 43|08|OW|1|Opacity Lookup Table Data
0029|WG12 Supplement 43|0b|SQ|1|Enhanced Palette Color Lookup Table Sequence
0029|WG12 Supplement 43|0c|SQ|1|Opacity 2 LUT Sequence
0029|WG12 Supplement 43|0d|CS|1|Opacity 2 LUT Transfer Function
0029|WG12 Supplement 43|0e|CS|1|Data Path ID
0029|WG12 Supplement 43|0f|CS|1|RGB LUT Transfer Function
0029|WG12 Supplement 43|10|CS|1|Alpha LUT Transfer Function
0041|WG12 Supplement 43|01|CS|1|Performed Protocol Type
0009|HMC - CT - ID|00|OB|1|Image ID Information Patient Name ID
0009|HMC - CT - ID|01|OB|1|Image ID Information Patient Comment
0019|SET WINDOW|00|SH|1|Set Window Image Filter
0019|SET WINDOW|01|US|1|Set Window Magnification Power
0017|SVISION|20|SQ|1|Scheduled Procedure Step List
0017|SVISION|a0|IS|1|Fixed Grid System
0017|SVISION|f0|IS|1|Images SOP Class
0019|SVISION|16|IS|1|Unknown
0019|SVISION|91|IS|1|Central Beam X
0019|SVISION|92|IS|1|Central Beam Y
0019|SVISION|93|IS|1|Tube Turn Angle
0019|SVISION|94|IS|1|Stand Drive Level
0019|SVISION|a0|DS|1|Extended Exposure Time
0019|SVISION|a1|DS|1|Actual Exposure Time
0019|SVISION|a8|DS|1|Extended X-ray Tube Current
0019|SVISION|b0|IS|1|Dose Indicator
0019|SVISION|b1|IS|1|Shift Reference Value
0019|SVISION|f0|IS|1|Unknown
0021|SVISION|50|DS|1|Minimal Window Latitude
0021|SVISION|51|DS|1|Maximal Window Latitude
0021|SVISION|52|DS|1|Relative Window Alignment
0021|SVISION|60|IS|1|Decomposition Layer
0023|SVISION|f0|IS|1|Image SOP Class
0025|SVISION|09|IS|1|Image Stitched Manually
0025|SVISION|0a|IS|1|Image Stitched Automatically
0029|SVISION|00|IS|1|Key Note Instance UID
0029|SVISION|01|IS|1|Storage State
0029|SVISION|02|IS|1|Referenced Image SOP Class
0029|SVISION|03|IS|1|Referenced Image Instance UID
0029|SVISION|04|IS|1|Related Presentation State Number
0029|SVISION|05|IS|1|Related Presentation State UID
5653|Vital Images SW 3.4|10|OB|1|Saved Workflow
5653|Vital Images SW 3.4|11|LO|1|Saved Workflow File Name
5653|Vital Images SW 3.4|12|OB|1|Saved Workflow File Data
5653|Vital Images SW 3.4|13|SL|1|Saved Workflow File Length
5653|Vital Images SW 3.4|14|SQ|1|Saved Workflow File Sequence
5653|Vital Images SW 3.4|15|SQ|1|Image Sequence
5653|Vital Images SW 3.4|16|SL|1|Volume Interpolated Slices
5653|Vital Images SW 3.4|17|UI|1|Volume SOP Instance UID
5653|Vital Images SW 3.4|18|SH|1|Saved Workflow Mark
5653|Vital Images SW 3.4|19|UI|1|Volume Study Instance UID
5653|Vital Images SW 3.4|20|SL|1|Number of Study Saved Workflow
5653|Vital Images SW 3.4|21|SL|1|Number of Series Saved Workflow
5653|Vital Images SW 3.4|22|UI|1|Volume Series Instance UID
5653|Vital Images SW 3.4|23|LO|1|Saved Workflow Code Meaning
5653|Vital Images SW 3.4|24|OB|1|Saved Workflow Data
5653|Vital Images SW 3.4|25|SL|1|Saved Workflow Data Length
0781|PI Private Block (0781:3000 - 0781:30FF)|01|US|1|Unknown
0781|PI Private Block (0781:3000 - 0781:30FF)|02|US|1|Unknown
0781|PI Private Block (0781:3000 - 0781:30FF)|05|FL|1|Unknown
0781|PI Private Block (0781:3000 - 0781:30FF)|09|FL|4|Unknown
0203|Riverain Medical|00|LO|1|Unknown
0203|Riverain Medical|01|LO|1|Unknown
0203|Riverain Medical|02|LO|1|Unknown
0203|Riverain Medical|03|LO|1|Unknown
0203|Riverain Medical|10|LO|1|Unknown
0203|Riverain Medical|f0|UI|1|Unknown
0203|Riverain Medical|f1|UI|1|Unknown
0029|INTELERAD MEDICAL SYSTEMS|16|US|1|Unknown
0029|INTELERAD MEDICAL SYSTEMS|17|US|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|01|LO|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|02|LO|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|03|UN|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|04|UN|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|05|UN|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|06|UN|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|07|UN|1|Unknown
0071|INTELERAD MEDICAL SYSTEMS INTELEVIEWER|0a|UN|1|Unknown
3f01|INTELERAD MEDICAL SYSTEMS|09|LO|1|Unknown
3f01|INTELERAD MEDICAL SYSTEMS|0a|DA|1|Unknown
3f01|INTELERAD MEDICAL SYSTEMS|0b|TM|1|Unknown
3f03|INTELERAD MEDICAL SYSTEMS|01|SQ|1|Unknown
3f03|INTELERAD MEDICAL SYSTEMS|02|DT|1|Unknown
3f03|INTELERAD MEDICAL SYSTEMS|03|LO|1|Unknown
3f03|INTELERAD MEDICAL SYSTEMS|04|LO|1|Unknown
4453|DR Systems, Inc.|00|LO|1|Exam ?
4453|DR Systems, Inc.|01|LO|1|Exam ID
4453|DR Systems, Inc.|02|LO|1|Image Type
4453|DR Systems, Inc.|04|LO|1|File Type
4453|DR Systems, Inc.|05|LO|1|File Suffix
4453|DR Systems, Inc.|0a|LO|1|Annotation Type
4453|DR Systems, Inc.|0c|SQ|1|Original Instance UID Sequence
0859|ETIAM DICOMDIR|40|DS|1|Unknown
0077|TERARECON AQUARIUS|10|UI|1-n|Original Series/Study UID
0077|TERARECON AQUARIUS|12|UI|1-n|Original SOP UID
0077|TERARECON AQUARIUS|14|LO|1-n|Referenced Volume ID
0077|TERARECON AQUARIUS|16|CS|1|Binary Data Name SCS
0077|TERARECON AQUARIUS|20|LO|1-n|Binary Data Name
0077|TERARECON AQUARIUS|22|CS|1-n|Number of SOP Instance UID
0077|TERARECON AQUARIUS|24|CS|1-n|Number of Series Instance UID
0077|TERARECON AQUARIUS|26|US|1|Number of Binary Data
0077|TERARECON AQUARIUS|28|CS|1-n|Binary Data Type
0077|TERARECON AQUARIUS|30|UL|1-n|Binary Data Size
0077|TERARECON AQUARIUS|32|LO|1-n|Binary Data SubType
0077|TERARECON AQUARIUS|40|LO|1-n|Additional Information
0077|TERARECON AQUARIUS|50|OB|1|First Binary Data
0077|TERARECON AQUARIUS|60|OB|1|First Thumbnail
0077|TERARECON AQUARIUS|70|LO|1|Algorithm ID
0077|TERARECON AQUARIUS|80|LO|1|Volume ID
0077|TERARECON AQUARIUS|84|LO|1-n|COF Object UID
0077|TERARECON AQUARIUS|86|LO|1-n|Workflow Scene Status
0077|TERARECON AQUARIUS|88|UI|1-n|Reference SOP Instance UIDs
0077|TERARECON AQUARIUS|90|FL|1|COF Refinement Level
0009|EMAGEON STUDY HOME|00|LO|1|Unknown
0009|EMAGEON STUDY HOME|01|LO|1|Unknown
0009|EMAGEON JPEG2K INFO|00|SQ|1|Unknown
0009|EMAGEON JPEG2K INFO|01|DT|1|Unknown
0029|RadWorksMarconi|24|US|1-n|Key Frame Indices
0009|MeVis eatDicom|10|LO|1|eatDicom Version
0009|MeVis eatDicom|11|ST|1|eatDicom Options
0021|MeVis eD: Timepoint Information|10|LT|1|Timepoint DateTime
0021|MeVis eD: Timepoint Information|11|CS|1|Timepoint DateTime Type
0021|MeVis eD: Timepoint Information|12|UN|1|Timepoint Series Description
0021|MeVis eD: Timepoint Information|13|UN|1|Timepoint Gradient Directions
0021|MeVis eD: Timepoint Information|71|UN|1|Timepoint Empty Frames
0021|MeVis eD: Absolute Temporal Positions|10|LT|1|Timepoint DateTime
0021|MeVis eD: Absolute Temporal Positions|11|CS|1|Timepoint DateTime Type
0021|MeVis eD: Absolute Temporal Positions|12|UN|1|Timepoint Series Description
0021|MeVis eD: Absolute Temporal Positions|13|UN|1|Timepoint Gradient Directions
0021|MeVis eD: Absolute Temporal Positions|71|UN|1|Timepoint Empty Frames
0021|MeVis eD: Geometry Information|10|UN|1|Geometry Scanner Origin
0021|MeVis eD: Slice Information|10|UI|1-n|Slice SOP Instance UIDs
0029|ShowcaseAppearance|10|DS|1|Unknown
0029|ShowcaseAppearance|11|DS|1|Unknown
0029|ShowcaseAppearance|12|DS|1|Unknown
0029|ShowcaseAppearance|13|DS|1|Unknown
0029|ShowcaseAppearance|14|SQ|1|Unknown
0099|NQHeader|01|UI|1|Version
0099|NQHeader|02|UI|1|Analyzed Series UID
0099|NQHeader|03|LT|1|License
0099|NQHeader|04|SS|1|Return Code
0099|NQHeader|05|LT|1|Return Message
0099|NQHeader|10|FL|1|MI
0099|NQHeader|20|SH|1|Units
0099|NQHeader|21|FL|1|ICV
0199|NQLeft|01|FL|1|Left Cortical White Matter
0199|NQLeft|02|FL|1|Left Cortical Gray Matter
0199|NQLeft|03|FL|1|Left 3rd Ventricle
0199|NQLeft|04|FL|1|Left 4th Ventricle
0199|NQLeft|05|FL|1|Left 5th Ventricle
0199|NQLeft|06|FL|1|Left Lateral Ventricle
0199|NQLeft|07|FL|1|Left Inferior Lateral Ventricle
0199|NQLeft|08|FL|1|Left Inferior CSF
0199|NQLeft|09|FL|1|Left Cerebellar White Matter
0199|NQLeft|0a|FL|1|Left Cerebellar Gray Matter
0199|NQLeft|0b|FL|1|Left Hippocampus
0199|NQLeft|0c|FL|1|Left Amygdala
0199|NQLeft|0d|FL|1|Left Thalamus
0199|NQLeft|0e|FL|1|Left Caudate
0199|NQLeft|0f|FL|1|Left Putamen
0199|NQLeft|10|FL|1|Left Pallidum
0199|NQLeft|11|FL|1|Left Ventral Diencephalon
0199|NQLeft|14|FL|1|Left Exterior CSF
0199|NQLeft|15|FL|1|Left WM Hypo
0199|NQLeft|16|FL|1|Left Other
0199|NQLeft|17|FL|1|Left Cortex Unkown
0199|NQLeft|18|FL|1|Left Cortex Bankssts
0199|NQLeft|19|FL|1|Left Cortex Caudal Anterior Cingulate
0199|NQLeft|1a|FL|1|Left Cortex Caudal Middle Frontal
0199|NQLeft|1b|FL|1|Left Cortex Corpus Callosum
0199|NQLeft|1c|FL|1|Left Cortex Cuneus
0199|NQLeft|1d|FL|1|Left Cortex Entorhinal
0199|NQLeft|1e|FL|1|Left Cortex Fusiform
0199|NQLeft|1f|FL|1|Left Cortex Inferior Parietal
0199|NQLeft|20|FL|1|Left Cortex Inferior Temporal
0199|NQLeft|21|FL|1|Left Cortex Isthmus Cingulate
0199|NQLeft|22|FL|1|Left Cortex Lateral Occipital
0199|NQLeft|23|FL|1|Left Cortex Lateral Orbito Frontal
0199|NQLeft|24|FL|1|Left Cortex Lingual
0199|NQLeft|25|FL|1|Left Cortex Medial Orbito Frontal
0199|NQLeft|26|FL|1|Left Cortex Middle Temporal
0199|NQLeft|27|FL|1|Left Cortex Parahippocampal
0199|NQLeft|28|FL|1|Left Cortex Paracentral
0199|NQLeft|29|FL|1|Left Cortex Pars Opercularis
0199|NQLeft|2a|FL|1|Left Cortex Pars Orbitalis
0199|NQLeft|2b|FL|1|Left Cortex Pars Triangularis
0199|NQLeft|2c|FL|1|Left Cortex Pericalcarine
0199|NQLeft|2d|FL|1|Left Cortex Postcentral
0199|NQLeft|2e|FL|1|Left Cortex Posterior Cingulate
0199|NQLeft|2f|FL|1|Left Cortex Precentral
0199|NQLeft|30|FL|1|Left Cortex Precuneus
0199|NQLeft|31|FL|1|Left Cortex Rostral Anterior Cingulate
0199|NQLeft|32|FL|1|Left Cortex Rostral Middle Frontal
0199|NQLeft|33|FL|1|Left Cortex Superior Frontal
0199|NQLeft|34|FL|1|Left Cortex Superior Parietal
0199|NQLeft|35|FL|1|Left Cortex Superior Temporal
0199|NQLeft|36|FL|1|Left Cortex Supramarginal
0199|NQLeft|37|FL|1|Left Cortex Frontal Pole
0199|NQLeft|38|FL|1|Left Cortex Temporal Pole
0199|NQLeft|39|FL|1|Left Cortex Transvere Temporal
0199|NQLeft|3a|FL|1|Left Meningie
0299|NQRight|01|FL|1|Right Cortical White Matter
0299|NQRight|02|FL|1|Right Cortical Gray Matter
0299|NQRight|03|FL|1|Right 3rd Ventricle
0299|NQRight|04|FL|1|Right 4th Ventricle
0299|NQRight|05|FL|1|Right 5th Ventricle
0299|NQRight|06|FL|1|Right Lateral Ventricle
0299|NQRight|07|FL|1|Right Inferior Lateral Ventricle
0299|NQRight|08|FL|1|Right Inferior CSF
0299|NQRight|09|FL|1|Right Cerebellar White Matter
0299|NQRight|0a|FL|1|Right Cerebellar Gray Matter
0299|NQRight|0b|FL|1|Right Hippocampus
0299|NQRight|0c|FL|1|Right Amygdala
0299|NQRight|0d|FL|1|Right Thalamus
0299|NQRight|0e|FL|1|Right Caudate
0299|NQRight|0f|FL|1|Right Putamen
0299|NQRight|10|FL|1|Right Pallidum
0299|NQRight|11|FL|1|Right Ventral Diencephalon
0299|NQRight|12|FL|1|Right Nucleus Accumbens
0299|NQRight|13|FL|1|Right Brain Stem
0299|NQRight|14|FL|1|Right Exterior CSF
0299|NQRight|15|FL|1|Right WM Hypo
0299|NQRight|16|FL|1|Right Other
0299|NQRight|17|FL|1|Right Cortex Unkown
0299|NQRight|18|FL|1|Right Cortex Bankssts
0299|NQRight|19|FL|1|Right Cortex Caudal Anterior Cingulate
0299|NQRight|1a|FL|1|Right Cortex Caudal Middle Frontal
0299|NQRight|1b|FL|1|Right Cortex Corpus Callosum
0299|NQRight|1c|FL|1|Right Cortex Cuneus
0299|NQRight|1d|FL|1|Right Cortex Entorhinal
0299|NQRight|1e|FL|1|Right Cortex Fusiform
0299|NQRight|1f|FL|1|Right Cortex Inferior Parietal
0299|NQRight|20|FL|1|Right Cortex Inferior Temporal
0299|NQRight|21|FL|1|Right Cortex Isthmus Cingulate
0299|NQRight|22|FL|1|Right Cortex Lateral Occipital
0299|NQRight|23|FL|1|Right Cortex Lateral Orbito Frontal
0299|NQRight|24|FL|1|Right Cortex Lingual
0299|NQRight|25|FL|1|Right Cortex Medial Orbito Frontal
0299|NQRight|26|FL|1|Right Cortex Middle Temporal
0299|NQRight|27|FL|1|Right Cortex Parahippocampal
0299|NQRight|28|FL|1|Right Cortex Paracentral
0299|NQRight|29|FL|1|Right Cortex Pars Opercularis
0299|NQRight|2a|FL|1|Right Cortex Pars Orbitalis
0299|NQRight|2b|FL|1|Right Cortex Pars Triangularis
0299|NQRight|2c|FL|1|Right Cortex Pericalcarine
0299|NQRight|2d|FL|1|Right Cortex Postcentral
0299|NQRight|2e|FL|1|Right Cortex Posterior Cingulate
0299|NQRight|2f|FL|1|Right Cortex Precentral
0299|NQRight|30|FL|1|Right Cortex Precuneus
0299|NQRight|31|FL|1|Right Cortex Rostral Anterior Cingulate
0299|NQRight|32|FL|1|Right Cortex Rostral Middle Frontal
0299|NQRight|33|FL|1|Right Cortex Superior Frontal
0299|NQRight|34|FL|1|Right Cortex Superior Parietal
0299|NQRight|35|FL|1|Right Cortex Superior Temporal
0299|NQRight|36|FL|1|Right Cortex Supramarginal
0299|NQRight|37|FL|1|Right Cortex Frontal Pole
0299|NQRight|38|FL|1|Right Cortex Temporal Pole
0299|NQRight|39|FL|1|Right Cortex Transvere Temporal
0299|NQRight|3a|FL|1|Right Meningie
0055|VEPRO VIF 3.0 DATA|20|OB|1|Unknown
0055|VEPRO VIF 3.0 DATA|30|OB|1|Icon Data
0055|VEPRO VIF 3.0 DATA|65|OB|1|Image Hash Value
0055|VEPRO VIM 5.0 DATA|10|OB|1|Unknown
0055|VEPRO VIM 5.0 DATA|20|OB|1|Unknown
0055|VEPRO VIM 5.0 DATA|30|OB|1|Icon Data
0055|VEPRO VIM 5.0 DATA|51|UI|1|Unknown
0055|VEPRO VIM 5.0 DATA|65|OB|1|Image Hash Value
0057|VEPRO BROKER 1.0|10|SQ|1|Data Replace Sequence
0057|VEPRO BROKER 1.0 DATA REPLACE|20|SQ|1|Original Data Sequence
0057|VEPRO BROKER 1.0 DATA REPLACE|30|SQ|1|Replaced Data Sequence
0057|VEPRO BROKER 1.0 DATA REPLACE|40|DA|1|Date of Data Replacement
0057|VEPRO BROKER 1.0 DATA REPLACE|41|TM|1|Time of Data Replacement
0057|VEPRO BROKER 1.0 DATA REPLACE|42|LO|1|Dicom Receive Node
0057|VEPRO BROKER 1.0 DATA REPLACE|43|LO|1|Application Name
0057|VEPRO BROKER 1.0 DATA REPLACE|44|LO|1|Computer Name
0059|VEPRO DICOM TRANSFER 1.0|10|SQ|1|Dicom Transfer Info
0059|VEPRO DICOM RECEIVE DATA 1.0|40|DA|1|Receive Date
0059|VEPRO DICOM RECEIVE DATA 1.0|41|TM|1|Receive Time
0031|KONICA1.0|49|UN|1|Unknown
0013|CTP|11|LO|1|Trial Name
0013|CTP|12|LO|1|Site Name
0013|CTP|13|LO|1|Site ID
0059|VEPRO DICOM RECEIVE DATA 1.0|42|ST|1|Receive Node
0059|VEPRO DICOM RECEIVE DATA 1.0|43|ST|1|Receive Application
0059|VEPRO DICOM RECEIVE DATA 1.0|50|ST|1|Receive Local Computer
0059|VEPRO DICOM RECEIVE DATA 1.0|51|ST|1|Receive Local AE Title
0059|VEPRO DICOM RECEIVE DATA 1.0|60|ST|1|Receive Remote Computer
0059|VEPRO DICOM RECEIVE DATA 1.0|61|ST|1|Receive Remote AE Title
0059|VEPRO DICOM RECEIVE DATA 1.0|70|UI|1|Receive Original Transfer Syntax
0043|dcm4che/archive|10|OB|1|Patient Pk
0043|dcm4che/archive|11|OB|1|Study Pk
0043|dcm4che/archive|12|OB|1|Series Pk
0043|dcm4che/archive|13|OB|1|Instance Pk
0043|dcm4che/archive|14|AE|1|Calling AE Title
0043|dcm4che/archive|15|AE|1|Called AE Title
0043|dcm4che/archive|16|DT|1|Instance Updated
0043|dcm4che/archive|20|SQ|1|Work Item Sequence
0043|dcm4che/archive|30|UI|1|Dcm4che URI Referenced Transfer Syntax UID
1269|IMS s.r.l. Biopsy Private Code|01|IS|1|Biopsy Image
1269|IMS s.r.l. Biopsy Private Code|10|IS|1-n|Biopsy Markers X
1269|IMS s.r.l. Biopsy Private Code|11|IS|1-n|Biopsy Markers Y
1269|IMS s.r.l. Biopsy Private Code|12|IS|1-n|Biopsy Markers Number
1269|IMS s.r.l. Biopsy Private Code|20|IS|1|Biopsy Area Left Border
1269|IMS s.r.l. Biopsy Private Code|21|IS|1|Biopsy Area Right Border
1269|IMS s.r.l. Biopsy Private Code|22|IS|1|Biopsy Area Top Border
1269|IMS s.r.l. Biopsy Private Code|23|IS|1|Biopsy Area Bottom Border
1269|IMS s.r.l. Biopsy Private Code|24|IS|1|Biopsy Number
1271|IMS s.r.l. Mammography Private Code|01|IS|1|Threshold 1
1271|IMS s.r.l. Mammography Private Code|02|IS|1|Threshold 2
1271|IMS s.r.l. Mammography Private Code|10|IS|1|Segmentation Left Border
1271|IMS s.r.l. Mammography Private Code|11|IS|1|Segmentation Right Border
1271|IMS s.r.l. Mammography Private Code|12|IS|1|Segmentation Top Border
1271|IMS s.r.l. Mammography Private Code|13|IS|1|Segmentation Bottom Border
1271|IMS s.r.l. Mammography Private Code|20|IS|1|Compressor Status
1271|IMS s.r.l. Mammography Private Code|21|IS|1|Collimator Type
1271|IMS s.r.l. Mammography Private Code|22|IS|1|Biopsy Specimen
1271|IMS s.r.l. Mammography Private Code|30|IS|1|Printer Segmentation
1271|IMS s.r.l. Mammography Private Code|31|IS|1|Printer 8x10 Format
1271|IMS s.r.l. Mammography Private Code|32|FD|1|Printer 8x10 Size X
1271|IMS s.r.l. Mammography Private Code|33|FD|1|Printer 8x10 Size Y
1271|IMS s.r.l. Mammography Private Code|34|IS|1|Printer 8x10 Area Left Border
1271|IMS s.r.l. Mammography Private Code|35|IS|1|Printer 8x10 Area Right Border
1271|IMS s.r.l. Mammography Private Code|36|IS|1|Printer 8x10 Area Top Border
1271|IMS s.r.l. Mammography Private Code|37|IS|1|Printer 8x10 Area Bottom Border
0031|KONICA1.0|4a|UN|1|Unknown
1271|IMS s.r.l. Mammography Private Code|38|LO|1|Rotation And Inclination Sensor Presence
1271|IMS s.r.l. Mammography Private Code|39|US|1-n|Window Center For For Processing Images
1271|IMS s.r.l. Mammography Private Code|40|US|1-n|Window Width For For Processing Images
1271|IMS s.r.l. Mammography Private Code|41|LO|1-n|Window Center and Width Explanation For For Processing Images
1271|IMS s.r.l. Mammography Private Code|42|LT|1|Processing Information
1271|IMS s.r.l. Mammography Private Code|43|LT|1|Filename
1271|IMS s.r.l. Mammography Private Code|44|LT|1|Contrast View
1271|IMS s.r.l. Mammography Private Code|45|IS|1|Threshold 3
1271|IMS s.r.l. Mammography Private Code|46|IS|1|Threshold 4
1271|IMS s.r.l. Mammography Private Code|47|IS|1|Threshold 5
1271|IMS s.r.l. Mammography Private Code|48|IS|1|Threshold 6
1271|IMS s.r.l. Mammography Private Code|49|IS|1|Threshold 7
1271|IMS s.r.l. Mammography Private Code|50|IS|1|Threshold 8
1271|IMS s.r.l. Mammography Private Code|51|IS|1|Threshold 9
1271|IMS s.r.l. Mammography Private Code|52|IS|1|Threshold 9
1271|IMS s.r.l. Mammography Private Code|53|IS|1|Scaling Factor For Processing
1271|IMS s.r.l. Mammography Private Code|54|IS|1|ConfirmX Image
1271|IMS s.r.l. Mammography Private Code|55|IS|1|Background counts
1271|IMS s.r.l. Mammography Private Code|56|IS|1|WL Roi Area X
1271|IMS s.r.l. Mammography Private Code|57|IS|1|WL Roi Area Y
1271|IMS s.r.l. Mammography Private Code|60|IS|1|Second Processing Image
1271|IMS s.r.l. Mammography Private Code|61|IS|1|S Filter
1271|IMS s.r.l. Mammography Private Code|62|IS|1|U Filter
1271|IMS s.r.l. Mammography Private Code|63|IS|1|Anonymous
1271|IMS s.r.l. Mammography Private Code|70|IS|1|Tomo SAD
1271|IMS s.r.l. Mammography Private Code|71|IS|1|Tomo Detector YAW
1271|IMS s.r.l. Mammography Private Code|72|IS|1|Tomo Detector Pitch
1271|IMS s.r.l. Mammography Private Code|73|IS|1|Tomo Detector Roll
1271|IMS s.r.l. Mammography Private Code|74|IS|1|Tomo Focal Spot X
1271|IMS s.r.l. Mammography Private Code|75|IS|1|Tomo Focal Spot Y
1271|IMS s.r.l. Mammography Private Code|76|IS|1|Tomo Xray Start Angle
1271|IMS s.r.l. Mammography Private Code|77|IS|1|Tomo Xray End Angle
1271|IMS s.r.l. Mammography Private Code|78|IS|1|Tomo Xray Angle
1271|IMS s.r.l. Mammography Private Code|79|IS|1|Tomo Exposure Counter
1271|IMS s.r.l. Mammography Private Code|80|IS|1|Tomo Exposure Number
1271|IMS s.r.l. Mammography Private Code|81|IS|1|Tomo WL Modified
1271|IMS s.r.l. Mammography Private Code|82|IS|1|Tomo Projection
1271|IMS s.r.l. Mammography Private Code|83|IS|1|Key Object Selection Title Code
0031|KONICA1.0|4b|UN|1|Unknown
1271|IMS s.r.l. Mammography Private Code|84|IS|1|Rejected for Quality Reasons Code
1271|IMS s.r.l. Mammography Private Code|85|IS|1|Unknown
0031|KONICA1.0|00|LO|1|Unknown
0031|KONICA1.0|01|US|1|Unknown
0031|KONICA1.0|05|US|1|Unknown
0031|KONICA1.0|06|LO|1|Unknown
0031|KONICA1.0|08|LO|1|Unknown
0031|KONICA1.0|09|US|1|Unknown
0031|KONICA1.0|0a|LO|1|Unknown
0031|KONICA1.0|0b|US|1|Unknown
0031|KONICA1.0|0c|US|1|Unknown
0031|KONICA1.0|0d|US|1|Unknown
0031|KONICA1.0|0e|US|1|Unknown
0031|KONICA1.0|10|US|1|Unknown
0031|KONICA1.0|11|US|1|Unknown
0031|KONICA1.0|12|US|1|Unknown
0031|KONICA1.0|13|US|1|Unknown
0031|KONICA1.0|14|US|1|Unknown
0031|KONICA1.0|15|US|1|Unknown
0031|KONICA1.0|16|US|1|Unknown
0031|KONICA1.0|17|US|1|Unknown
0031|KONICA1.0|18|US|1|Unknown
0031|KONICA1.0|19|US|1|Unknown
0031|KONICA1.0|1a|US|1|Unknown
0031|KONICA1.0|1b|US|1|Unknown
0031|KONICA1.0|1c|US|1|Unknown
0031|KONICA1.0|1d|US|1|Unknown
0031|KONICA1.0|1e|LO|1|Unknown
0031|KONICA1.0|20|SQ|1|Unknown
0031|KONICA1.0|21|SQ|1|Unknown
0031|KONICA1.0|22|SQ|1|Unknown
0031|KONICA1.0|23|SQ|1|Unknown
0031|KONICA1.0|24|SQ|1|Unknown
0031|KONICA1.0|25|SQ|1|Unknown
0031|KONICA1.0|26|SQ|1|Unknown
0031|KONICA1.0|27|SQ|1|Unknown
0031|KONICA1.0|28|SQ|1|Unknown
0031|KONICA1.0|29|SQ|1|Unknown
0031|KONICA1.0|2a|SQ|1|Unknown
0031|KONICA1.0|2b|SQ|1|Unknown
0031|KONICA1.0|2c|SQ|1|Unknown
0031|KONICA1.0|2d|SQ|1|Unknown
0031|KONICA1.0|2e|SQ|1|Unknown
0031|KONICA1.0|2f|SQ|1|Unknown
0031|KONICA1.0|30|US|1|Unknown
0031|KONICA1.0|31|US|1|Unknown
0031|KONICA1.0|32|US|1|Unknown
0031|KONICA1.0|33|US|1|Unknown
0031|KONICA1.0|34|US|1|Unknown
0031|KONICA1.0|35|UN|1|Unknown
0031|KONICA1.0|36|UN|1|Unknown
0031|KONICA1.0|37|US|1|Unknown
0031|KONICA1.0|38|US|1|Unknown
0031|KONICA1.0|39|US|1|Unknown
0031|KONICA1.0|3a|UN|1|Unknown
0031|KONICA1.0|3b|US|1|Unknown
0031|KONICA1.0|3c|US|1|Unknown
0031|KONICA1.0|3d|US|1|Unknown
0031|KONICA1.0|3e|US|1|Unknown
0031|KONICA1.0|3f|US|1|Unknown
0031|KONICA1.0|40|US|1|Unknown
0031|KONICA1.0|41|US|1|Unknown
0031|KONICA1.0|42|US|1|Unknown
0031|KONICA1.0|44|US|1|Unknown
0031|KONICA1.0|45|US|1|Unknown
0031|KONICA1.0|46|US|1|Unknown
0031|KONICA1.0|47|US|1|Unknown
0031|KONICA1.0|48|US|1|Unknown
0031|KONICA1.0|4c|UN|1|Unknown
0031|KONICA1.0|4d|US|1|Unknown
0031|KONICA1.0|4e|US|1|Unknown
0031|KONICA1.0|4f|US|1|Unknown
0031|KONICA1.0|50|US|1|Unknown
0031|KONICA1.0|51|US|1|Unknown
0031|KONICA1.0|52|US|1|Unknown
0031|KONICA1.0|53|US|1|Unknown
0031|KONICA1.0|54|US|1|Unknown
0031|KONICA1.0|55|US|1|Unknown
0031|KONICA1.0|56|UN|1|Unknown
0031|KONICA1.0|57|US|1|Unknown
0031|KONICA1.0|58|US|1|Unknown
0031|KONICA1.0|59|US|1|Unknown
0031|KONICA1.0|5a|US|1|Unknown
0031|KONICA1.0|5b|US|1|Unknown
0031|KONICA1.0|5c|UN|1|Unknown
0031|KONICA1.0|62|US|1|Unknown
0031|KONICA1.0|63|US|3|Unknown
0031|KONICA1.0|6b|US|1|Unknown
0031|KONICA1.0|70|US|1|Unknown
0031|KONICA1.0|71|LO|1|Unknown
0031|KONICA1.0|72|US|1|Unknown
0031|KONICA1.0|73|UN|1|Unknown
0031|KONICA1.0|74|LO|1|Unknown
0031|KONICA1.0|75|UN|1|Unknown
0031|KONICA1.0|77|UN|1|Unknown
0031|KONICA1.0|78|UN|1|Unknown
0031|KONICA1.0|79|UN|1|Unknown
0031|KONICA1.0|7a|UN|1|Unknown
0031|KONICA1.0|7b|UN|1|Unknown
0031|KONICA1.0|7c|UN|1|Unknown
0031|KONICA1.0|7d|UN|1|Unknown
0031|KONICA1.0|7e|UN|1|Unknown
0031|KONICA1.0|7f|UN|1|Unknown
0031|KONICA1.0|80|UN|1|Unknown
0031|KONICA1.0|81|UN|1|Unknown
0031|KONICA1.0|82|UN|1|Unknown
0031|KONICA1.0|83|UN|1|Unknown
0031|KONICA1.0|84|UN|1|Unknown
0031|KONICA1.0|85|UN|1|Unknown
0031|KONICA1.0|86|UN|1|Unknown
0031|KONICA1.0|87|UN|1|Unknown
0031|KONICA1.0|88|UN|1|Unknown
0031|KONICA1.0|89|UN|1|Unknown
0031|KONICA1.0|8a|UN|1|Unknown
0031|KONICA1.0|8b|UN|1|Unknown
0031|KONICA1.0|8c|US|1|Unknown
0031|KONICA1.0|8d|US|1|Unknown
0031|KONICA1.0|8e|LO|1|Unknown
0031|KONICA1.0|8f|UN|1|Unknown
0031|KONICA1.0|90|UN|1|Unknown
0031|KONICA1.0|91|US|1|Unknown
0031|KONICA1.0|92|UN|1|Unknown
0031|KONICA1.0|93|UN|1|Unknown
0031|KONICA1.0|94|UN|1|Unknown
0031|KONICA1.0|95|UN|1|Unknown
0031|KONICA1.0|a1|IS|2|Unknown
0031|KONICA1.0|a2|IS|1|Unknown
0031|KONICA1.0|a5|US|1|Unknown
0031|KONICA1.0|a6|US|1|Unknown
0031|KONICA1.0|a7|UN|1|Unknown
0031|KONICA1.0|a8|US|1|Unknown
0031|KONICA1.0|aa|US|1|Unknown
0031|KONICA1.0|ab|DA|1|Unknown
0031|KONICA1.0|ac|TM|1|Unknown
0031|KONICA1.0|ad|DA|1|Unknown
0031|KONICA1.0|ae|TM|1|Unknown
0031|KONICA1.0|b0|US|1|Unknown
0031|KONICA1.0|b1|US|1|Unknown
0031|KONICA1.0|b2|US|1|Unknown
0031|KONICA1.0|b3|US|1|Unknown
0031|KONICA1.0|b4|US|1|Unknown
0031|KONICA1.0|b5|US|1|Unknown
0031|KONICA1.0|b6|US|1|Unknown
0031|KONICA1.0|b7|UN|1|Unknown
0031|KONICA1.0|b8|LO|1|Unknown
0031|KONICA1.0|b9|LO|1|Unknown
0031|KONICA1.0|ba|US|1|Unknown
0031|KONICA1.0|bc|US|1|Unknown
0031|KONICA1.0|be|UN|1|Unknown
0031|KONICA1.0|bf|US|1|Unknown
0031|KONICA1.0|c0|UN|1|Unknown
0031|KONICA1.0|c1|UN|1|Unknown
0031|KONICA1.0|c2|UN|1|Unknown
0031|KONICA1.0|c3|UN|1|Unknown
0031|KONICA1.0|c4|UN|1|Unknown
0031|KONICA1.0|c5|UN|1|Unknown
0031|KONICA1.0|c6|UN|1|Unknown
0031|KONICA1.0|c7|UN|1|Unknown
0031|KONICA1.0|c8|UN|1|Unknown
0031|KONICA1.0|c9|UN|1|Unknown
0031|KONICA1.0|ca|UN|1|Unknown
0031|KONICA1.0|cb|UN|1|Unknown
0031|KONICA1.0|cc|UN|1|Unknown
0031|KONICA1.0|cd|UN|1|Unknown
0031|KONICA1.0|ce|US|1|Unknown
0031|KONICA1.0|cf|US|1|Unknown
0031|KONICA1.0|d0|UN|1|Unknown
0031|KONICA1.0|d1|UN|1|Unknown
0031|KONICA1.0|d2|UN|1|Unknown
0031|KONICA1.0|d3|UN|1|Unknown
0031|KONICA1.0|d4|US|1|Unknown
0031|KONICA1.0|d5|UN|1|Unknown
0031|KONICA1.0|d6|UN|1|Unknown
0031|KONICA1.0|d7|US|1|Unknown
0031|KONICA1.0|d8|US|1|Unknown
0031|KONICA1.0|d9|LO|1|Unknown
0031|KONICA1.0|da|UN|1|Unknown
0031|KONICA1.0|db|UN|1|Unknown
0031|KONICA1.0|dc|UN|1|Unknown
0031|KONICA1.0|dd|UN|1|Unknown
0031|KONICA1.0|de|UN|1|Unknown
0031|KONICA1.0|df|UN|1|Unknown
0031|KONICA1.0|e0|UN|1|Unknown
0031|KONICA1.0|e1|US|1|Unknown
0031|KONICA1.0|e2|UN|1|Unknown
0031|KONICA1.0|e3|UN|1|Unknown
0031|KONICA1.0|e4|UN|1|Unknown
0031|KONICA1.0|e5|US|1|Unknown
0031|KONICA1.0|e6|UN|1|Unknown
0031|KONICA1.0|f0|US|1|Unknown
0031|KONICA1.0|ff|SQ|1|Private Data Sequence
0009|DZDICOM 4.3.0|01|UI|1|Unknown
0009|DZDICOM 4.3.0|02|LO|1|Unknown
0009|DZDICOM 4.3.0|03|LO|1|Unknown
0009|DZDICOM 4.3.0|04|IS|1|Unknown
0009|DZDICOM 4.3.0|05|LO|1|Unknown
0009|DZDICOM 4.3.0|06|LO|1|Unknown
0009|DZDICOM 4.3.0|07|LO|1|Unknown
0009|DZDICOM 4.3.0|08|IS|1|Unknown
0009|DZDICOM 4.3.0|11|LO|1|Unknown
0009|DZDICOM 4.3.0|12|LO|1|Unknown
0009|DZDICOM 4.3.0|13|LO|1|Unknown
0009|DZDICOM 4.3.0|14|LO|1|Unknown
0009|DZDICOM 4.3.0|15|LO|1|Unknown
0009|DZDICOM 4.3.0|16|LO|1|Unknown
0009|DZDICOM 4.3.0|17|LO|1|Unknown
0009|DZDICOM 4.3.0|70|IS|1|Unknown
0009|DZDICOM 4.3.0|71|IS|1|Unknown
0009|DZDICOM 4.3.0|72|IS|1|Unknown
0009|DZDICOM 4.3.0|74|IS|1|Unknown
0009|DZDICOM 4.3.0|7a|IS|1|Unknown
0009|DZDICOM 4.3.0|a1|LO|1|Unknown
0009|DZDICOM 4.3.0|a2|IS|1|Unknown
0009|DZDICOM 4.3.0|f1|LO|1|Unknown
0009|DZDICOM 4.3.0|f7|IS|1|Unknown
0009|DZDICOM 4.3.0|f9|IS|1|Unknown
0019|FOEM 1.0|50|IS|1|Unknown
0025|FOEM 1.0|10|US|1|Unknown
0025|FOEM 1.0|12|US|1|Unknown
0029|FOEM 1.0|20|IS|1|Unknown
5533|Visus Change|33|SQ|1|Save Sequence
5533|Visus Change|35|DA|1|Save Date
5533|Visus Change|37|LO|1|Save Originator
5533|Visus Change|39|FD|1|Save ID
5533|Visus Change|3b|TM|1|Save Time
0099|SYNARC_1.0|01|OB|1|Unknown
0099|SYNARC_1.0|02|OB|1|Unknown
0099|SYNARC_1.0|03|LO|1|Unknown
0099|SYNARC_1.0|04|US|1-n|Unknown
0099|SYNARC_1.0|05|LO|1|Unknown
0011|PixelMed Publishing|02|UC|1|Strain Description
0011|PixelMed Publishing|03|LO|1|Strain Nomenclature
0011|PixelMed Publishing|04|LO|1|Strain Stock Number
0011|PixelMed Publishing|05|SQ|1|Strain Source Registry Code Sequence
0011|PixelMed Publishing|06|SQ|1|Strain Stock Sequence
0011|PixelMed Publishing|07|LO|1|Strain Source
0011|PixelMed Publishing|08|UT|1|Strain Additional Information
0011|PixelMed Publishing|20|SQ|1|Strain Code Sequence
0011|PixelMed Publishing|50|LO|1|Cell Line Designation
0011|PixelMed Publishing|51|SQ|1|Cell Line Tissue of Origin Code Sequence
0011|PixelMed Publishing|52|SQ|1|Cell Line Histologic Type Code Sequence
0011|PixelMed Publishing|53|SQ|1|Cell Line Species of Origin Code Sequence
0011|PixelMed Publishing|54|UL|1|Cell Line Number of Passages
0011|PixelMed Publishing|71|SQ|1|Source Patient Group Identification Sequence
0011|PixelMed Publishing|72|SQ|1|Group of Patients Identification Sequence
0011|PixelMed Publishing|73|US|3|Subject Relative Position in Image
0021|PixelMed Publishing|01|SQ|1|Unassigned Shared Converted Attributes Sequence
0021|PixelMed Publishing|02|SQ|1|Unassigned Per-Frame Converted Attributes Sequence
0021|PixelMed Publishing|03|SQ|1|Conversion Source Attributes Sequence
0041|PixelMed Publishing|01|SQ|1|Quantity Definition Code Sequence
7fe1|PixelMed Publishing|01|OF|1|Float Pixel Data
7fe1|PixelMed Publishing|02|OD|1|Double Pixel Data
0011|METAEMOTION GINKGO|01|LT|1|KeyFile Indicator
0011|METAEMOTION GINKGO|0b|LT|1|Serialized Diagnose and Markers
0011|METAEMOTION GINKGO RETINAL|01|LT|1|KeyFile Indicator
0011|METAEMOTION GINKGO RETINAL|0b|LT|1|Serialized Diagnose and Markers
0011|METAEMOTION GINKGO RETINAL|0c|UN|1|Virtual Aneritra Contrast Image
0055|PMOD_1|01|FD|1-n|Frame Start Times Vector
0055|PMOD_1|02|FD|3-3n|Frame Positions Vector
0055|PMOD_1|03|FD|6-6n|Frame Orientations Vector
0055|PMOD_1|04|FD|1-n|Frame Durations Vector
0055|PMOD_1|05|FD|1-n|Frame Rescale Slope Vector
7fe1|PMOD_GENPET|01|UT|1|Slices Names
7fe1|PMOD_GENPET|02|UT|1|Gene Codes
7fe1|PMOD_GENPET|03|UT|1|Gene Labels
0011|ULTRAVISUAL_TAG_SET1|01|CS|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|02|UN|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|03|UN|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|08|LO|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|10|US|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|11|UN|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|12|UI|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|18|UL|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|19|UN|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|1a|CS|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|1b|IS|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|1c|IS|1|Unknown
0011|ULTRAVISUAL_TAG_SET1|1d|LO|1|Unknown
0015|MATAKINA_10|28|LO|1|Volpara Density Grade
0015|MATAKINA_10|29|LT|1|Volpara Run Information
0015|MATAKINA_10|30|LO|1|Volpara Density Grade Cutoffs
0101|PM|05|LO|1-n|Image Enhancement Parameter File
0101|PM|06|IS|1|Original Sigmoid Ratio
0863|Biospace Med : EOS Tag|10|SL|1|Image Type
0863|Biospace Med : EOS Tag|23|SL|1|Calibration Flag
0863|Biospace Med : EOS Tag|26|UL|1|Attribute Version
0863|Biospace Med : EOS Tag|27|SL|1|Resizing Flag
0863|Biospace Med : EOS Tag|28|SL|1|Logarithm Flag
0863|Biospace Med : EOS Tag|32|SL|1|Left Collimator Edge
0863|Biospace Med : EOS Tag|33|SL|1|Right Collimator Edge
0863|Biospace Med : EOS Tag|34|FL|1|Distance Source to Patient of Biplane Pair
0863|Biospace Med : EOS Tag|35|SL|1|Line Correction Flag
0863|Biospace Med : EOS Tag|36|SL|1|Contrast Enhancement Flag
0863|Biospace Med : EOS Tag|37|SL|1|Calibre Value
0863|Biospace Med : EOS Tag|38|SL|1|High Frequency Line Correction Max Threshold
0863|Biospace Med : EOS Tag|39|SL|1|High Frequency Line Correction Min Threshold
0863|Biospace Med : EOS Tag|40|FL|1|Greater Limit
0863|Biospace Med : EOS Tag|41|FL|1|Lower Limit
0863|Biospace Med : EOS Tag|42|FL|1|Frontal Detector Blades Opening
0863|Biospace Med : EOS Tag|43|FL|1|Frontal Tube Blades Opening
0863|Biospace Med : EOS Tag|44|FL|1|Lateral Detector Blades Opening
0863|Biospace Med : EOS Tag|45|FL|1|Lateral Tube Blades Opening
0863|Biospace Med : EOS Tag|46|DS|1-n|ThreeD Calibration Parameters
0863|Biospace Med : EOS Tag|57|CS|1|Image Horizontal Flip
0019|PRIVATE_CODE_STRING_0019|00|FD|1|Calibration
0019|PRIVATE_CODE_STRING_0019|01|FD|1|Depth Conversion
0019|PRIVATE_CODE_STRING_0019|02|FD|1|Stepsize
0019|PRIVATE_CODE_STRING_0019|03|SL|1-n|Warning
0019|PRIVATE_CODE_STRING_0019|04|ST|1|DataID
0021|PRIVATE_CODE_STRING_0021|70|FD|1|Distance Base Plane to Template
0021|PRIVATE_CODE_STRING_0021|71|FD|16|Volume to Patient Matrix
0021|PRIVATE_CODE_STRING_0021|72|FD|16|Patient to World Matrix
0021|PRIVATE_CODE_STRING_0021|73|SL|1|Base Plane
0021|PRIVATE_CODE_STRING_0021|74|SL|1|Reference Plane
0021|PRIVATE_CODE_STRING_0021|75|SL|1|Apex Plane
0021|PRIVATE_CODE_STRING_0021|76|FD|1|Base Plane Offset
1001|PRIVATE_CODE_STRING_1001|a0|SQ|1|Marker Sequence
1001|PRIVATE_CODE_STRING_1001|a1|SL|1|Marker Type
1001|PRIVATE_CODE_STRING_1001|a2|SL|1|Marker Number
1001|PRIVATE_CODE_STRING_1001|a3|FD|3|Marker 3D Position
1001|PRIVATE_CODE_STRING_1001|b0|SL|1|Distance Unit
1001|PRIVATE_CODE_STRING_1001|b1|SL|1|Dose Unit
1001|PRIVATE_CODE_STRING_1001|b2|SL|1|Normalisation Mode
1001|PRIVATE_CODE_STRING_1001|b3|FD|1|Normalisation Factor
1001|PRIVATE_CODE_STRING_1001|b4|FD|1|F-Value
1001|PRIVATE_CODE_STRING_1001|b5|FD|1|Prescribed Dose
1001|PRIVATE_CODE_STRING_1001|b6|FD|1|Absolute Dose Factor
1001|PRIVATE_CODE_STRING_1001|b7|SL|1|Decoupled sk
1001|PRIVATE_CODE_STRING_1001|b8|FD|1|Absolute Time Factor
1001|PRIVATE_CODE_STRING_1001|b9|FD|1|Total Treatment Time
1001|PRIVATE_CODE_STRING_1001|ba|SL|1|TG 43 Model
1001|PRIVATE_CODE_STRING_1001|bb|SL|1|3D Dose Grid Size
1001|PRIVATE_CODE_STRING_1001|bc|FD|3|Dose Grid Corner 1
1001|PRIVATE_CODE_STRING_1001|bd|FD|3|Dose Grid Corner 2
1001|PRIVATE_CODE_STRING_1001|be|FD|1|Patient Data Conversion
1001|PRIVATE_CODE_STRING_1001|bf|FD|1|Volume Data Conversion
1001|PRIVATE_CODE_STRING_1001|c0|FD|3|Volume Data Vector
1001|PRIVATE_CODE_STRING_1001|c1|SL|1|Optimization Method
1001|PRIVATE_CODE_STRING_1001|c2|SL|1|Display Method
1001|PRIVATE_CODE_STRING_1001|c3|SL|1|Geometrical Method
1001|PRIVATE_CODE_STRING_1001|c5|SL|1|VOI Number
1001|PRIVATE_CODE_STRING_1001|c6|LO|1|VOI Name
1001|PRIVATE_CODE_STRING_1001|c7|SL|1|VOI Type
1001|PRIVATE_CODE_STRING_1001|c8|SL|1|VOI Class
1001|PRIVATE_CODE_STRING_1001|c9|SL|1|VOI Priority
1001|PRIVATE_CODE_STRING_1001|ca|SL|1|No of Points
1001|PRIVATE_CODE_STRING_1001|cb|FD|1|Percent On Surface
1001|PRIVATE_CODE_STRING_1001|cc|FD|1|Surface Margin
1001|PRIVATE_CODE_STRING_1001|cd|SL|1|Selected
1001|PRIVATE_CODE_STRING_1001|ce|FD|1|Dose Limit
1001|PRIVATE_CODE_STRING_1001|cf|FD|1|Importance Factor
1001|PRIVATE_CODE_STRING_1001|d0|FD|1|Importance Factor From
1001|PRIVATE_CODE_STRING_1001|d1|FD|1|Importance Factor To
1001|PRIVATE_CODE_STRING_1001|d2|FD|1|Focus
1001|PRIVATE_CODE_STRING_1001|d3|SL|1|Surface Sampling Method
1001|PRIVATE_CODE_STRING_1001|d4|FD|1|Number of Sampling Points Per ccm
1001|PRIVATE_CODE_STRING_1001|d5|SL|1|Convergence Accuracy
3335|CAD Sciences|07|UN|1|Unknown
1001|PRIVATE_CODE_STRING_1001|d6|SL|1|Max No of Convergence Iterations
1001|PRIVATE_CODE_STRING_1001|d7|FD|1|Weight Smoothing
1001|PRIVATE_CODE_STRING_1001|d8|SL|1|Steps Per Importance Factor
1001|PRIVATE_CODE_STRING_1001|d9|FD|1|Constraints PTVDmax
1001|PRIVATE_CODE_STRING_1001|da|FD|1|Constraints NTDmax
1001|PRIVATE_CODE_STRING_1001|db|SL|1|Algorithmic Population Size
1001|PRIVATE_CODE_STRING_1001|dc|SL|1|Algorithmic Generations
1001|PRIVATE_CODE_STRING_1001|dd|SL|1|Algorithmic Initializations
1001|PRIVATE_CODE_STRING_1001|de|SL|1|Min No Of SDP
1001|PRIVATE_CODE_STRING_1001|df|SL|1|Depth Method
1001|PRIVATE_CODE_STRING_1001|e0|SL|1|Depth Defined On
1001|PRIVATE_CODE_STRING_1001|e1|FD|1|Depth
1001|PRIVATE_CODE_STRING_1001|e2|SQ|1|VOI Based Placement Settings Sequence
1001|PRIVATE_CODE_STRING_1001|e7|SL|1|VOI Selected
1001|PRIVATE_CODE_STRING_1001|e8|FD|1|Margin
1001|PRIVATE_CODE_STRING_1001|e9|SL|1|Selection Method
1001|PRIVATE_CODE_STRING_1001|ea|FD|1|Selection Distance
1001|PRIVATE_CODE_STRING_1001|eb|FD|1|WBT On Contour Spacing
1001|PRIVATE_CODE_STRING_1001|ec|FD|1|WBT Urethra Margin
1001|PRIVATE_CODE_STRING_1001|ed|FD|1|WBT Searching Radius PTV
1001|PRIVATE_CODE_STRING_1001|ee|FD|1|WBT Searching Radius OAR
1001|PRIVATE_CODE_STRING_1001|ef|FD|3|WBT Starting Point
1001|PRIVATE_CODE_STRING_1001|f0|FD|4|WBT Surface
1001|PRIVATE_CODE_STRING_1001|f1|FD|4|WBT No of Interior Catheters
1001|PRIVATE_CODE_STRING_1001|f2|FD|4|WBT Relative Radius
1001|PRIVATE_CODE_STRING_1001|f3|SL|1|Sorting Method
1003|PRIVATE_CODE_STRING_1003|01|UN|1|Number Of Probes
1003|PRIVATE_CODE_STRING_1003|10|UN|1|US Probe Sequence
1003|PRIVATE_CODE_STRING_1003|11|UN|1|Identifier
1003|PRIVATE_CODE_STRING_1003|12|UN|1|Probe Name
1003|PRIVATE_CODE_STRING_1003|13|UN|1|Depth
1003|PRIVATE_CODE_STRING_1003|14|UN|1|Frequency
1003|PRIVATE_CODE_STRING_1003|15|UN|1|Gain
1003|PRIVATE_CODE_STRING_1003|16|UN|1|Power
1003|PRIVATE_CODE_STRING_1003|17|UN|1|Dynamic Range
1003|PRIVATE_CODE_STRING_1003|18|UN|1|Frame Averaging
1003|PRIVATE_CODE_STRING_1003|19|UN|1|Field Of View
1003|PRIVATE_CODE_STRING_1003|20|UN|1|TGC
1003|PRIVATE_CODE_STRING_1003|2a|UN|1|Number Of Focus Sets
1003|PRIVATE_CODE_STRING_1003|2b|UN|1|Current Focus Set
1003|PRIVATE_CODE_STRING_1003|2c|UN|1|Image Enhancement Filter Index
1003|PRIVATE_CODE_STRING_1003|2d|UN|1|Rejection Filter Low
1003|PRIVATE_CODE_STRING_1003|2e|UN|1|Rejection Filter High
1003|PRIVATE_CODE_STRING_1003|2f|UN|1|Brightness
1003|PRIVATE_CODE_STRING_1003|30|UN|1|Contrast
1003|PRIVATE_CODE_STRING_1003|31|UN|1|Gamma
1003|PRIVATE_CODE_STRING_1003|32|UN|1|Speckle Enabled
1003|PRIVATE_CODE_STRING_1003|33|UN|1|Speckle Level
1003|PRIVATE_CODE_STRING_1003|40|UN|1|Focus Set Sequence
1003|PRIVATE_CODE_STRING_1003|41|UN|1|Identifier
1003|PRIVATE_CODE_STRING_1003|42|UN|1|Number Of Focus Zone
1003|PRIVATE_CODE_STRING_1003|43|UN|1|Focus
3007|PRIVATE_CODE_STRING_3007|00|FD|16|Volume to Patient Matrix
3007|PRIVATE_CODE_STRING_3007|01|FD|16|Volume Resolution Conversion
3007|PRIVATE_CODE_STRING_3007|02|FD|16|Volume Data Conversion
3007|PRIVATE_CODE_STRING_3007|03|FD|16|Patient Data Conversion
3007|PRIVATE_CODE_STRING_3007|04|FD|16|DICOM Data Conversion
300b|PRIVATE_CODE_STRING_300B|00|SL|1|Template Mode
300b|PRIVATE_CODE_STRING_300B|01|LO|1|Template ID
300b|PRIVATE_CODE_STRING_300B|02|SL|1|Number of Columns
300b|PRIVATE_CODE_STRING_300B|03|FD|1|Column Distance
300b|PRIVATE_CODE_STRING_300B|04|SL|1|Number of Rows
300b|PRIVATE_CODE_STRING_300B|05|FD|1|Row Distance
300b|PRIVATE_CODE_STRING_300B|06|SL|1|Origin
300b|PRIVATE_CODE_STRING_300B|07|SH|1-n|Column Numbering
300b|PRIVATE_CODE_STRING_300B|08|SH|1-n|Row Numbering
300b|PRIVATE_CODE_STRING_300B|09|SS|1-n|Used Holes Array
300b|PRIVATE_CODE_STRING_300B|0a|SL|1|Lock Status
300b|PRIVATE_CODE_STRING_300B|0c|UN|1|Identifier
300b|PRIVATE_CODE_STRING_300B|0d|UN|1|Modification Type
300b|PRIVATE_CODE_STRING_300B|0e|UN|1|Modification Value
300b|PRIVATE_CODE_STRING_300B|0f|UN|1|Transformation Matrix
000d|INSTRU_PRIVATE_IDENT_CODE|00|OB|1|Image Xml Data
000d|SCANORA_PRIVATE_IDENT_CODE|00|OB|1|Image Xml Data
0019|NNT|02|US|1|Unknown
0019|NNT|03|DS|1|Unknown
0019|NNT|04|DS|1|Unknown
0019|NNT|05|DS|1|Unknown
0019|NNT|06|DS|1|Unknown
0019|NNT|07|DS|1|Unknown
0019|NNT|09|DS|1|Unknown
0019|NNT|0a|DS|1|Unknown
0019|NNT|0b|DS|1|Unknown
0019|NNT|0c|DS|1|Unknown
0019|NNT|0d|DS|1|Unknown
0019|NNT|0e|DS|1|Unknown
0019|NNT|0f|DS|1|Unknown
0019|NNT|12|DS|1|Unknown
0019|NNT|13|DS|1|Unknown
0019|NNT|1e|DS|3|Unknown
0019|NNT|1f|DS|1|Unknown
0019|NNT|20|DS|1|Unknown
0019|NNT|21|DS|1|Unknown
0019|NNT|22|IS|1|Unknown
0019|NNT|23|IS|1|Unknown
0019|NNT|24|LO|1|Unknown
0019|NNT|25|IS|1|Unknown
0019|NNT|26|LO|1|Unknown
0019|NNT|27|LO|1|Unknown
0019|NNT|28|LO|1|Unknown
0019|NNT|30|LO|1|Unknown
0019|NNT|31|IS|1|Unknown
0019|NNT|32|IS|1|Unknown
0019|NNT|33|DS|8|Unknown
3335|CAD Sciences|00|UN|1|Unknown
3335|CAD Sciences|06|UN|1|Unknown
3335|CAD Sciences|08|UN|1|Unknown
3335|iCAD PK|10|LO|1|Unknown
3335|iCAD PK|15|LO|1|Unknown
3335|iCAD PK|16|LO|1|Unknown
3335|iCAD PK|17|LO|1|Unknown
3335|iCAD PK|18|LO|1|Unknown
3335|iCAD PK|2a|LO|1|Unknown
3335|iCAD PK|34|LO|1|Unknown
3335|iCAD PK|35|LO|1|Unknown
3335|iCAD PK|3b|LO|1|Unknown
3335|iCAD PK|40|LO|1|Unknown
3335|iCAD PK|50|LO|1|Unknown
3335|iCAD PK|51|LO|1|Unknown
3335|iCAD PK|52|LO|1|Unknown
3335|iCAD PK|53|LO|1|Unknown
3335|iCAD PK|54|LO|1|Unknown
3335|iCAD PK|55|LO|1|Unknown
3335|iCAD PK|56|LO|1|Unknown
3335|iCAD PK|57|LO|1|Unknown
3335|iCAD PK|70|LO|1|Unknown
3335|iCAD PK|71|LO|1|Unknown
3335|iCAD PK|72|LO|1|Unknown
3335|iCAD PK|73|LO|1|Unknown
3335|iCAD PK|74|LO|1|Unknown
3335|iCAD PK|75|UN|1|Unknown
3335|iCAD PK|80|LO|1|Unknown
3335|iCAD PK|81|LO|1|Unknown
3335|iCAD PK|82|LO|1|Unknown
3335|iCAD PK|83|LO|1|Unknown
3335|iCAD PK|84|LO|1|Unknown
3335|iCAD PK|85|LO|1|Unknown
3335|iCAD PK|86|LO|1|Unknown
3335|iCAD PK|87|LO|1|Unknown
3335|iCAD PK|88|LO|1|Unknown
3335|iCAD PK|89|LO|1|Unknown
3335|iCAD PK|8a|LO|1|Unknown
3335|iCAD PK|8b|LO|1|Unknown
3335|iCAD PK|8c|LO|1|Unknown
3335|iCAD PK|8d|LO|1|Unknown
3335|iCAD PK|8e|LO|1|Unknown
3335|iCAD PK|8f|LO|1|Unknown
3335|iCAD PK|90|LO|1|Unknown
3335|iCAD PK|91|LO|1|Unknown
3335|iCAD PK|92|LO|1|Unknown
3335|iCAD PK|93|LO|1|Unknown
3335|iCAD PK|94|LO|1|Unknown
3335|iCAD PK|95|LO|1|Unknown
3335|iCAD PK|a0|LO|1|Unknown
3335|iCAD PK|a1|LO|1|Unknown
3335|iCAD PK|a2|LO|1|Unknown
3335|iCAD PK|a3|LO|1|Unknown
3335|iCAD PK|a4|LO|1|Unknown
3335|iCAD PK|a5|LO|1|Unknown
3335|iCAD PK|a6|LO|1|Unknown
3335|iCAD PK|a7|LO|1|Unknown
3335|iCAD PK|a8|LO|1|Unknown
3335|iCAD PK|a9|LO|1|Unknown
3335|iCAD PK|aa|LO|1|Unknown
3335|iCAD PK|ab|LO|1|Unknown
3335|iCAD PK|ac|LO|1|Unknown
3335|iCAD PK|ad|LO|1|Unknown
3335|iCAD PK|ae|LO|1|Unknown
3335|iCAD PK|af|LO|1|Unknown
3335|iCAD PK|b0|LO|1|Unknown
3335|iCAD PK|b1|LO|1|Unknown
3335|iCAD PK|c0|LO|1|Unknown
3335|iCAD PK Study|00|LO|1|Unknown
3335|iCAD PK Study|01|LO|1|Unknown
3335|iCAD PK Study|02|LO|1|Unknown
3335|iCAD PK Study|03|LO|1|Unknown
3335|iCAD PK Study|04|LO|1|Unknown
3335|iCAD PK Study|05|LO|1|Unknown
3335|iCAD PK Study|06|LO|1|Unknown
3335|iCAD PK Study|07|LO|1|Unknown
3335|iCAD PK Study|08|LO|1|Unknown
3335|iCAD PK Study|09|LO|1|Unknown
3335|iCAD PK Study|0a|LO|1|Unknown
3335|iCAD PK Study|0b|LO|1|Unknown
3335|iCAD PK Study|0c|LO|1|Unknown
3335|iCAD PK Study|0d|LO|1|Unknown
3335|iCAD PK Study|0e|LO|1|Unknown
3335|iCAD PK Study|0f|LO|1|Unknown
3335|iCAD PK Study|10|LO|1|Unknown
3335|iCAD PK Study|11|LO|1|Unknown
3335|iCAD PK Study|12|LO|1|Unknown
3335|iCAD PK Study|13|LO|1|Unknown
3335|iCAD PK Study|14|LO|1|Unknown
3335|iCAD PK Study|15|LO|1|Unknown
3335|iCAD PK Study|16|LO|1|Unknown
3335|iCAD PK Study|17|LO|1|Unknown
3335|iCAD PK Study|18|LO|1|Unknown
3335|iCAD PK Study|19|LO|1|Unknown
3335|iCAD PK Study|1a|LO|1|Unknown
3335|iCAD PK Study|1b|LO|1|Unknown
7fdf|TomTec|50|OB|1|Unknown
7fdf|TomTec|51|OB|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|15|LO|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|16|LO|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|17|LO|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|18|UT|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|19|IS|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|1a|IS|1|Unknown
0029|CARESTREAM IMAGE INFORMATION|1b|IS|1|Unknown
ffff|Carestream Health TIFF|ff|UN|1|Unknown
3111|RamSoft File Kind Identifier|10|CS|1|Binary Document Type
3113|RamSoft Custom Report Identifier|10|OB|1|Binary Document
3113|RamSoft Custom Report Identifier|20|UL|1|Binary Document Size
3129|RamSoft Race Identifier|10|LO|1|Unknown
0011|MDDX|01|UT|1|AES Encrypted Values
0011|MDDX|02|LO|1|Allup Version Details
0011|MDDX|03|LO|1|Mask Id
7fe1|MDDX|01|UT|1|AES Encrypted Values
7fe1|MDDX|02|LO|1|Allup Version Details
7fe1|MDDX|03|LO|1|Mask Id
0099|QTUltrasound|00|SS|1|Breast Density Value
0009|BioscanMedisoScivisNanoSPECT|35|DS|1|Unknown
0009|MEDISO-1|30|DT|1|Unknown
0009|MEDISO-1|36|FD|1|Unknown
0009|MEDISO-1|c0|FD|1|Unknown
0009|MEDISO-1|c1|OB|1|Unknown
0009|MEDISO-1|c4|OB|1|Unknown
0009|MEDISO-1|d2|LO|1|Unknown
0009|MEDISO-1|d5|LO|1|Unknown
0009|MEDISO-1|dc|SQ|1|Unknown
0009|MEDISO-1|de|UL|1|Unknown
0009|MEDISO-1|df|UL|1|Unknown
0009|MEDISO-1|e0|US|1|Unknown
0009|MEDISO-1|e1|FD|1|Unknown
0009|MEDISO-1|e6|OB|1|Unknown
0009|MEDISO-1|e9|UI|1-n|Unknown
0009|MEDISO-1|ee|DT|1|Unknown
0009|MEDISO-1|ef|DT|1|Unknown
0009|MEDISO-1|f0|FD|1|Unknown
0009|MEDISO-1|f1|FD|1|Unknown
0009|MEDISO-1|f2|FD|1|Unknown
0009|MEDISO-1|f3|FD|1|Unknown
0009|MEDISO-1|fa|ST|1|Unknown
0009|MEDISO-1|fb|US|1|Unknown
0011|MEDISO-1|06|LO|1|Unknown
6001|SCIVIS-1|a0|DS|1|Unknown
6001|SCIVIS-1|a1|DS|1|Unknown
6001|SCIVIS-1|a2|US|1|Unknown
6001|SCIVIS-1|a3|DS|1|Unknown
6001|SCIVIS-1|a4|IS|1|Unknown
6001|SCIVIS-1|a5|ST|1|Unknown
6001|SCIVIS-1|a6|ST|1|Unknown
6001|SCIVIS-1|a7|FL|1|Unknown
6001|SCIVIS-1|a8|FL|1|Unknown
6001|SCIVIS-1|a9|IS|1|Unknown
6001|SCIVIS-1|aa|IS|1|Unknown
6001|SCIVIS-1|ab|ST|1|Unknown
0009|Brainlab-S9-History|31|SQ|1|Unknown
0009|Brainlab-S9-History|32|SQ|1|Unknown
0009|Brainlab-S9-History|33|SQ|1|Unknown
0063|Brainlab-S32-SO|01|LO|1|Unknown
0063|Brainlab-S32-SO|10|SQ|1|Unknown
0073|Brainlab-S23-ProjectiveFusion|10|SQ|1|Projective Registration Sequence
0009|SPI Release 1|08|CS|1|Unknown
0009|PHILIPS MR/PART 12|2110|US|1|Unknown
0009|SPI-P Release 1|10|LO|1|Unknown
0009|SPI-P Release 1|a0|UN|1|Unknown
0011|SPI-P Release 1|20|UN|1|Unknown
0011|SPI-P Release 1|30|UN|1|Unknown
0019|PHILIPS MR/PART 7|00|IS|1|Unknown
0019|SPI-P-CTBE Release 1|00|IS|1|Unknown
0019|SPI-P-Private-DiDi Release 1|00|LT|1|Post Mode String
0019|SPI-P-XSB-VISUB Release 1|00|UN|1|Unknown
0019|PHILIPS MR/PART|1001|DS|1|Unknown
0019|SPI-P-Private-DiDi Release 1|01|LT|1|Post Data
0019|PHILIPS MR/PART|1002|DS|1|Unknown
0019|SPI-P-CTBE Release 1|02|IS|1|Unknown
0019|PHILIPS MR/PART|1003|DS|1|Unknown
0019|SPI-P-CTBE Release 1|03|DS|1|Unknown
0019|SPI-P-CTBE Release 1|04|IS|1|Unknown
0019|SPI-P-CTBE Release 1|05|DS|1|Unknown
0019|SPI-P-CTBE Release 1|0b|DS|1|Unknown
0019|SPI-P-CTBE Release 1|0c|IS|1|Unknown
0019|PHILIPS MR/PART 6|10|IS|1|Unknown
0019|SPI-P-PCR Release 2|10|US|1|Unknown
0019|SPI-P-Private-DiDi Release 1|10|LT|1|Image Header
0019|SPI-P-XSB-VISUB Release 1|10|UN|1|Unknown
0019|SPI-P-XSB-VISUB Release 1|11|UN|1|Unknown
0019|SPI-P-XSB-VISUB Release 1|12|UN|1|Unknown
0019|PHILIPS MR/PART|1014|CS|1|Unknown
0019|SPI-P-CTBE Release 1|14|IS|1|Unknown
0019|SPI-P-CTBE Release 1|18|IS|1|Unknown
0019|SPI-P-CTBE Release 1|19|IS|1|Unknown
0019|SPI-P-CTBE Release 1|1a|DS|1|Unknown
0019|SPI-P-CTBE Release 1|1b|IS|1|Unknown
0019|PHILIPS MR/PART|101c|CS|1|Unknown
0019|SPI-P-CTBE Release 1|1c|IS|1|Unknown
0019|PHILIPS MR/PART|101d|CS|1|Unknown
0019|SPI-P-CTBE Release 1|1d|DS|1|Unknown
0019|PHILIPS MR/PART|101e|DS|1|Unknown
0019|SPI-P-PCR Release 2|20|IS|1|Unknown
0019|SPI-P-XSB-VISUB Release 1|20|LO|1|Unknown
0019|PHILIPS MR/PART|1121|DS|1|Unknown
0019|SPI-P-PCR Release 2|21|LO|1|Unknown
0019|PHILIPS MR/PART|1123|DS|1-n|Unknown
0019|PHILIPS MR/PART|1124|DS|1-n|Unknown
0019|PHILIPS MR/PART|1125|DS|1-n|Unknown
0019|PHILIPS MR/PART|1126|DS|1-n|Unknown
0019|PHILIPS MR/PART|1127|DS|1-n|Unknown
0019|PHILIPS MR/PART|1128|CS|1|Unknown
0019|PHILIPS MR/PART|1129|DS|1-n|Unknown
0019|PHILIPS MR/PART|1130|LO|1-n|Unknown
0019|PHILIPS MR/PART|1131|DS|1-n|Unknown
0019|PHILIPS MR/PART|1040|US|1|Unknown
0019|SPI-P-PCR Release 2|40|DS|1|Unknown
0019|SPI-P-XSB-VISUB Release 1|40|UN|1|Unknown
0019|PHILIPS MR/PART|1050|IS|1|Unknown
0019|PHILIPS MR/PART|1150|DS|1|Unknown
0019|SPI-P-XSB-VISUB Release 1|50|LO|1|Unknown
0019|PHILIPS MR/PART|1151|DS|1|Unknown
0019|PHILIPS MR/PART|1152|DS|1|Unknown
0019|PHILIPS MR/PART|1153|IS|1|Unknown
0019|PHILIPS MR/PART|1154|DS|1|Unknown
0019|PHILIPS MR/PART|1155|DS|1|Unknown
0019|PHILIPS MR/PART|1156|DS|1|Unknown
0019|PHILIPS MR/PART|1157|US|1|Unknown
0019|PHILIPS MR/PART|1158|DS|1|Unknown
0019|PHILIPS MR/PART|1159|US|1|Unknown
0019|PHILIPS MR/PART|1160|DS|1|Unknown
0019|SPI-P-PCR Release 2|60|LO|1|Unknown
0019|PHILIPS MR/PART|1161|DS|1|Unknown
0019|PHILIPS MR/PART|1162|DS|1|Unknown
0019|PHILIPS MR/PART|1163|DS|1|Unknown
0019|PHILIPS MR/PART|1164|IS|1|Unknown
0019|PHILIPS MR/PART|1166|US|1|Unknown
0019|PHILIPS MR/PART|1067|US|1|Unknown
0019|PHILIPS MR/PART|1070|DS|1-n|Unknown
0019|SPI-P-PCR Release 2|80|US|1|Unknown
0019|DIDI TO PCR 1.1|89|IS|1|Exposure Index
0019|DIDI TO PCR 1.1|8a|IS|1|Collimator X
0019|PHILIPS MR/PART|108a|CS|1|Unknown
0019|DIDI TO PCR 1.1|8b|IS|1|Collimator Y
0019|PHILIPS MR/PART|108b|CS|1|Unknown
0019|DIDI TO PCR 1.1|8c|LO|1|Print Marker
0019|PHILIPS MR/PART|108c|CS|1|Unknown
0019|DIDI TO PCR 1.1|8d|LO|1|RGDV Name
0019|PHILIPS MR/PART|108d|CS|1|Unknown
0019|DIDI TO PCR 1.1|8e|LO|1|Acqd Sensitivity
0019|PHILIPS MR/PART|108e|CS|1|Unknown
0019|DIDI TO PCR 1.1|8f|LO|1|Processing Category
0019|PHILIPS MR/PART|108f|CS|1|Unknown
0019|SPI-P-PCR Release 2|90|LO|1|Unknown
0019|DIDI TO PCR 1.1|a0|LO|1|Version
0019|DIDI TO PCR 1.1|a1|LO|1|Ranging Mode
0019|DIDI TO PCR 1.1|a2|DS|1|Abdomen Brightness
0019|DIDI TO PCR 1.1|a3|DS|1|Fixed Brightness
0019|DIDI TO PCR 1.1|a4|DS|1|Detail Contrast
0019|DIDI TO PCR 1.1|a5|DS|1|Contrast Balance
0019|DIDI TO PCR 1.1|a6|DS|1|Structure Boost
0019|DIDI TO PCR 1.1|a7|DS|1|Structure Preference
0019|DIDI TO PCR 1.1|a8|DS|1|Noise Robustness
0019|DIDI TO PCR 1.1|a9|DS|1|Noise Dose Limit
0019|DIDI TO PCR 1.1|aa|DS|1|Noise Dose Step
0019|DIDI TO PCR 1.1|ab|DS|1|Noise Frequency Limit
0019|DIDI TO PCR 1.1|ac|DS|1|Weak Contrast Limit
0019|DIDI TO PCR 1.1|ad|DS|1|Strong Contrast Limit
0019|DIDI TO PCR 1.1|ae|DS|1|Structure Boost Offset
0019|DIDI TO PCR 1.1|af|LO|1|Smooth Gain
0019|DIDI TO PCR 1.1|b0|LO|1|Measure Field 1
0019|DIDI TO PCR 1.1|b1|LO|1|Measure Field 2
0019|DIDI TO PCR 1.1|b2|IS|1|Key Percentile 1
0019|DIDI TO PCR 1.1|b3|IS|1|Key Percentile 2
0019|DIDI TO PCR 1.1|b4|IS|1|Density LUT
0019|PHILIPS MR/PART|10b4|DS|1|Unknown
0019|DIDI TO PCR 1.1|b5|DS|1|Brightness
0019|PHILIPS MR/PART|10b5|DS|1|Unknown
0019|DIDI TO PCR 1.1|b6|DS|1|Gamma
0019|PHILIPS MR/PART|10b6|DS|1|Unknown
0019|PHILIPS MR/LAST|b7|IS|1|Unknown
0019|PHILIPS MR/PART|10d1|US|1|Unknown
0019|PHILIPS MR/PART|10d3|DS|1|Unknown
0019|PHILIPS MR/LAST|e4|IS|1|Unknown
0019|PHILIPS MR/LAST|e5|DS|1|Unknown
0019|PHILIPS MR/PART|10f0|IS|1|Unknown
0019|PHILIPS MR/PART|10f6|CS|1|Unknown
0019|PHILIPS MR/PART|10f7|CS|1|Unknown
0019|PHILIPS MR/PART|10f8|CS|1|Unknown
0019|PHILIPS MR/PART|10f9|CS|1|Unknown
0019|PHILIPS MR/PART|10fa|CS|1|Unknown
0019|PHILIPS MR/PART|10fb|CS|1|Unknown
0019|PHILIPS MR/PART|10fc|CS|1|Unknown
0019|SPI-P-PCR Release 2|a1|ST|1|Unknown
0019|SPI-P-PCR Release 2|a3|DS|1|Unknown
0019|SPI-P-PCR Release 2|a4|DS|1|Unknown
0019|SPI-P-PCR Release 2|a5|DS|1|Unknown
0019|SPI-P-PCR Release 2|a6|DS|1|Unknown
0019|SPI-P-PCR Release 2|a7|DS|1|Unknown
0019|SPI-P-PCR Release 2|a8|DS|1|Unknown
0019|SPI-P-PCR Release 2|a9|DS|1|Unknown
0019|SPI-P-PCR Release 2|aa|DS|1|Unknown
0019|SPI-P-PCR Release 2|ab|DS|1|Unknown
0019|SPI-P-PCR Release 2|ac|DS|1|Unknown
0019|SPI-P-PCR Release 2|ad|DS|1|Unknown
0019|SPI-P-PCR Release 2|ae|DS|1|Unknown
0019|SPI-P-PCR Release 2|af|ST|1|Unknown
0019|SPI-P-PCR Release 2|b0|ST|1|Unknown
0019|SPI-P-PCR Release 2|b1|ST|1|Unknown
0019|SPI-P-PCR Release 2|b2|IS|1|Unknown
0019|SPI-P-PCR Release 2|b3|IS|1|Unknown
0019|SPI-P-PCR Release 2|b4|IS|1|Unknown
0019|SPI-P-PCR Release 2|b5|DS|1|Unknown
0019|SPI-P-PCR Release 2|b6|DS|1|Unknown
0019|SPI-P-PCR Release 2|b7|ST|1|Unknown
0019|SPI-P-PCR Release 2|b8|DS|1|Unknown
0019|SPI-P-PCR Release 2|b9|ST|1|Unknown
0019|SPI-P-PCR Release 2|ba|ST|1|Unknown
0021|SPI-P-CTBE-Private Release 1|00|DS|1|Unknown
0021|PHILIPS MR/PART|1006|LO|1|Unknown
0021|PHILIPS MR/PART|1008|LO|1|Unknown
0021|PHILIPS MR/PART|1009|CS|1|Unknown
0021|PHILIPS MR/PART|100a|CS|1|Unknown
0021|PHILIPS MR/PART|100f|LO|1|Unknown
0021|PHILIPS MR/PART|1013|CS|1|Unknown
0021|PHILIPS MR/PART|1015|US|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|00|ST|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|00|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1;3|01|ST|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|01|DS|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|02|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1|0d|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|0e|SQ|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|0f|CS|1|Unknown
0029|SPI-P-Private_CDS Release 1|10|OB|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|10|LO|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|11|DS|1|Unknown
0029|SPI-P-Private_ICS Release 1|12|SQ|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|12|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1|1d|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|1e|SQ|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|1f|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1|20|UN|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|20|LO|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|21|DS|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|22|CS|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|2f|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|30|LT|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|30|LO|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|31|DS|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|32|CS|1|Unknown
0029|SPI-P-XSB-VISUB Release 1|3f|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1|4c|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|4d|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1|4e|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1|4f|FD|1|Unknown
0029|PHILIPS MR/PART|1050|DS|1|Unknown
0029|SPI-P-Private_ICS Release 1|50|FD|1|Unknown
0029|PHILIPS MR/PART|1051|DS|1|Unknown
0029|SPI-P-Private_ICS Release 1|51|FD|1|Unknown
0029|PHILIPS MR/PART|1052|DS|1|Unknown
0029|PHILIPS MR/PART|1053|DS|1|Unknown
0029|PHILIPS MR/LAST|62|IS|1|Unknown
0029|SPI-P-Private_ICS Release 1|6a|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1|6b|US|1|Unknown
0029|SPI-P-Private_ICS Release 1|72|SQ|1|Unknown
0029|SPI-P Release 1|90|DS|1-n|Unknown
0029|SPI-P Release 1|91|US|1|Unknown
0029|SPI-P-Private_ICS Release 1|91|IS|1|Unknown
0029|SPI-P Release 1|9f|CS|1|Unknown
0029|SPI-P Release 1|a0|DS|1-n|Unknown
0029|SPI-P-Private_ICS Release 1;2|a0|SL|1|Unknown
0029|SPI-P Release 1|a1|US|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|a1|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|a2|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|a3|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|a5|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|a6|SL|1|Unknown
0029|SPI-P Release 1|af|CS|1|Unknown
0029|SPI-P Release 1|b0|DS|1-n|Unknown
0029|SPI-P Release 1|b1|US|1|Unknown
0029|SPI-P Release 1|bf|CS|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|c0|SL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|c1|US|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|cb|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|cc|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|cd|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d0|UN|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d1|LO|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d2|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d3|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d4|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d5|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;1|d6|ST|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|d6|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|d7|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|d8|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;2|d9|SQ|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|d9|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|da|FL|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|dc|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|dd|FD|1|Unknown
0029|SPI-P-Private_ICS Release 1;4|e0|SQ|1|Unknown
0041|PHILIPS MR/LAST|07|LO|1|Unknown
0041|PHILIPS MR/LAST|09|DS|1|Unknown
0089|PMS-THORA-5.1|20|SQ|1|Unknown
0511|Philips PET Private Group|00|US|1|Private Data
0511|Philips PET Private Group|01|US|1|Private Data
0511|Philips PET Private Group|02|OB|1|Private Data
0511|Philips PET Private Group|03|OB|1|Private Data
0511|Philips PET Private Group|32|DS|1|Private Data
0511|Philips PET Private Group|50|DS|1|Private Data
1001|Philips Imaging DD 124|03|LO|1|Unknown
2001|Philips Imaging DD 129|00|SQ|1|Presentation State Sequence
2001|Philips Imaging DD 002|01|US|1|Unknown
2001|Philips Imaging DD 129|01|SQ|1|PresentationStateSequence
2001|Philips Imaging DD 002|02|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|05|SS|1|Graphic Annotation ParentID
2001|Philips Imaging DD 001|05|SS|1|Graphic Annotation ParentID
2001|PHILIPS IMAGING DD 001|09|FL|1|Image Prepulse Delay
2001|PHILIPS IMAGING DD 001|0c|CS|1|Arrhythmia Rejection
2001|PHILIPS IMAGING DD 001|0e|CS|1|Cardiac Cycled
2001|PHILIPS IMAGING DD 001|0f|SS|1|Cardiac Gate Width
2001|PHILIPS IMAGING DD 001|10|CS|1|Cardiac Sync
2001|Philips Imaging DD 002|13|SS|1|Unknown
2001|Philips Imaging DD 002|14|FD|1|Unknown
2001|Philips Imaging DD 002|15|FD|1|Unknown
2001|Philips Imaging DD 002|16|FD|1|Unknown
2001|Philips Imaging DD 002|17|FD|1|Unknown
2001|Philips Imaging DD 002|18|CS|1|Unknown
2001|Philips Imaging DD 002|19|FD|1|Unknown
2001|Philips Imaging DD 002|1a|FD|1|Unknown
2001|Philips Imaging DD 002|1b|FD|1|Unknown
2001|Philips Imaging DD 002|1c|FD|1|Unknown
2001|Philips Imaging DD 002|1d|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|1e|CS|1|Reformat Accuracy
2001|Philips Imaging DD 001|1e|CS|1|Reformat Accuracy
2001|Philips Imaging DD 002|1e|FD|1|Unknown
2001|Philips Imaging DD 002|1f|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|20|LO|1|Scanning Technique
2001|Philips Imaging DD 002|20|FD|1|Unknown
2001|Philips Imaging DD 002|21|FD|1|Unknown
2001|Philips Imaging DD 002|22|FD|1|Unknown
2001|Philips Imaging DD 002|23|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|24|CS|1|Series is Interactive
2001|Philips Imaging DD 002|24|FD|1|Unknown
2001|Philips Imaging DD 002|25|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|26|CS|1|Presentation State Subtraction Active
2001|Philips Imaging DD 001|26|CS|1|Presentation State Subtraction Active
2001|Philips Imaging DD 002|26|FD|1|Unknown
2001|Philips Imaging DD 001|20|LO|1|Scanning Technique
2001|Philips Imaging DD 001|24|CS|1|Series is Interactive
2001|Philips Imaging DD 002|27|FD|1|Unknown
2001|Philips Imaging DD 002|28|US|1|Unknown
2001|PHILIPS IMAGING DD 001|29|FL|1|Unknown
2001|Philips Imaging DD 001|29|FL|1|Unknown
2001|Philips Imaging DD 002|29|US|1|Unknown
2001|Philips Imaging DD 002|2a|US|1|Unknown
2001|PHILIPS IMAGING DD 001|2b|CS|1|Unknown
2001|Philips Imaging DD 001|2b|CS|1|Unknown
2001|Philips Imaging DD 002|2b|SS|1|Unknown
2001|Philips Imaging DD 002|2c|FD|1|Unknown
2001|Philips Imaging DD 002|2d|FD|1|Unknown
2001|Philips Imaging DD 002|2e|SS|1|Unknown
2001|Philips Imaging DD 002|2f|SS|1|Unknown
2001|Philips Imaging DD 002|30|SS|1|Unknown
2001|Philips Imaging DD 002|31|SS|1|Unknown
2001|Philips Imaging DD 002|32|SS|1|Unknown
2001|Philips Imaging DD 002|33|SS|1|Unknown
2001|Philips Imaging DD 002|34|SS|1|Unknown
2001|Philips Imaging DD 002|35|FD|1|Unknown
2001|Philips Imaging DD 002|36|FD|1|Unknown
2001|Philips Imaging DD 002|37|FD|1|Unknown
2001|PHILIPS IMAGING DD 001|39|FL|1|Unknown
2001|Philips Imaging DD 001|39|FL|1|Unknown
2001|Philips Imaging DD 002|39|CS|1|Unknown
2001|Philips Imaging DD 002|3a|SQ|1|Unknown
2001|Philips Imaging DD 002|3b|SQ|1|Unknown
2001|Philips Imaging DD 002|3c|SQ|1|Unknown
2001|PHILIPS IMAGING DD 001|3d|UL|1|Contour Fill Color
2001|Philips Imaging DD 001|3d|UL|1|Contour Fill Color
2001|Philips Imaging DD 002|3d|SQ|1|Unknown
2001|Philips Imaging DD 002|3e|SS|1|Unknown
2001|Philips Imaging DD 002|3f|SS|1|Unknown
2001|Philips Imaging DD 002|40|SS|1|Unknown
2001|PHILIPS IMAGING DD 001|43|IS|2|Ellipse Display Shutter Major Axis First End Point
2001|Philips Imaging DD 001|43|IS|2|Ellipse Display Shutter Major Axis First End Point
2001|PHILIPS IMAGING DD 001|44|IS|2|Ellipse Display Shutter Major Axis Second End Point
2001|Philips Imaging DD 001|44|IS|2|Ellipse Display Shutter Major Axis Second End Point
2001|PHILIPS IMAGING DD 001|45|IS|2|Ellipse Display Shutter Other Axis First End Point
2001|Philips Imaging DD 001|45|IS|2|Ellipse Display Shutter Other Axis First End Point
2001|PHILIPS IMAGING DD 001|46|CS|1|Graphic Line Style
2001|Philips Imaging DD 001|46|CS|1|Graphic Line Style
2001|PHILIPS IMAGING DD 001|47|FL|1|Graphic Line Width
2001|Philips Imaging DD 001|47|FL|1|Graphic Line Width
2001|PHILIPS IMAGING DD 001|48|SS|1|Graphic Annotation ID
2001|Philips Imaging DD 001|48|SS|1|Graphic Annotation ID
2001|PHILIPS IMAGING DD 001|4b|CS|1|Interpolation Method
2001|Philips Imaging DD 001|4b|CS|1|Interpolation Method
2001|PHILIPS IMAGING DD 001|4c|CS|1|Poly Line Begin Point Style
2001|Philips Imaging DD 001|4c|CS|1|Poly Line Begin Point Style
2001|PHILIPS IMAGING DD 001|4d|CS|1|Poly Line End Point Style
2001|Philips Imaging DD 001|4d|CS|1|Poly Line End Point Style
2001|PHILIPS IMAGING DD 001|4e|CS|1|Window Smoothing Taste
2001|Philips Imaging DD 001|4e|CS|1|Window Smoothing Taste
2001|PHILIPS IMAGING DD 001|50|LO|1|Graphic Marker Type
2001|Philips Imaging DD 001|50|LO|1|Graphic Marker Type
2001|PHILIPS IMAGING DD 001|51|IS|1|Overlay Plane ID
2001|Philips Imaging DD 001|51|IS|1|Overlay Plane ID
2001|PHILIPS IMAGING DD 001|52|UI|1|Image Presentation State UID
2001|Philips Imaging DD 001|52|UI|1|Image Presentation State UID
2001|PHILIPS IMAGING DD 001|53|CS|1|Presentation GL Transform Invert
2001|Philips Imaging DD 001|53|CS|1|Presentation GL Transform Invert
2001|PHILIPS IMAGING DD 001|54|FL|1|Contour Fill Transparency
2001|Philips Imaging DD 001|54|FL|1|Contour Fill Transparency
2001|PHILIPS IMAGING DD 001|55|UL|1|Graphic Line Color
2001|Philips Imaging DD 001|55|UL|1|Graphic Line Color
2001|PHILIPS IMAGING DD 001|56|CS|1|Graphic Type
2001|Philips Imaging DD 001|56|CS|1|Graphic Type
2001|PHILIPS IMAGING DD 001|58|UL|1|Contrast Transfer Taste
2001|PHILIPS IMAGING DD 001|5a|ST|1|Graphic Annotation Model
2001|Philips Imaging DD 001|5a|ST|1|Graphic Annotation Model
2001|PHILIPS IMAGING DD 001|5d|ST|1|Measurement Text Units
2001|Philips Imaging DD 001|5d|ST|1|Measurement Text Units
2001|PHILIPS IMAGING DD 001|5e|ST|1|Measurement Text Type
2001|Philips Imaging DD 001|5e|ST|1|Measurement Text Type
2001|PHILIPS IMAGING DD 001|64|SH|1|Text Type
2001|Philips Imaging DD 001|64|SH|1|Text Type
2001|PHILIPS IMAGING DD 001|65|SQ|1|Graphic Overlay Plane
2001|Philips Imaging DD 001|65|SQ|1|Graphic Overlay Plane
2001|PHILIPS IMAGING DD 001|67|CS|1|Linear Presentation GL Transform Shape Sub
2001|Philips Imaging DD 001|67|CS|1|Linear Presentation GL Transform Shape Sub
2001|PHILIPS IMAGING DD 001|68|SQ|1|Linear Modality GL Transform
2001|Philips Imaging DD 001|68|SQ|1|Linear Modality GL Transform
2001|PHILIPS IMAGING DD 001|69|SQ|1|Display Shutter
2001|Philips Imaging DD 001|69|SQ|1|Display Shutter
2001|PHILIPS IMAGING DD 001|6a|SQ|1|Spatial Transformation
2001|Philips Imaging DD 001|6a|SQ|1|Spatial Transformation
2001|PHILIPS IMAGING DD 001|6b|SQ|1|Unknown
2001|Philips Imaging DD 001|6b|SQ|1|Unknown
2001|PHILIPS IMAGING DD 001|6d|LO|1|Text Font
2001|Philips Imaging DD 001|6d|LO|1|Text Font
2001|PHILIPS IMAGING DD 001|6e|SH|1|Series Type
2001|Philips Imaging DD 001|6e|SH|1|Series Type
2001|PHILIPS IMAGING DD 001|71|CS|1|Graphic Constraint
2001|Philips Imaging DD 001|71|CS|1|Graphic Constraint
2001|PHILIPS IMAGING DD 001|72|IS|1|Ellipse Display Shutter Other Axis Second End Point
2001|Philips Imaging DD 001|72|IS|1|Ellipse Display Shutter Other Axis Second End Point
2001|Philips Imaging DD 002|72|FL|2|Unknown
2001|Philips Imaging DD 002|73|FL|2|Unknown
2001|PHILIPS IMAGING DD 001|74|DS|1|Unknown
2001|Philips Imaging DD 001|74|DS|1|Unknown
2001|PHILIPS IMAGING DD 001|75|DS|1|Unknown
2001|Philips Imaging DD 001|75|DS|1|Unknown
2001|PHILIPS IMAGING DD 001|76|UL|1|Number of Frames
2001|Philips Imaging DD 001|76|UL|1|Number of Frames
2001|PHILIPS IMAGING DD 001|77|CS|1|GL Transform Type
2001|Philips Imaging DD 001|77|CS|1|GL Transform Type
2001|PHILIPS IMAGING DD 001|7a|FL|1|Window Rounding Factor
2001|Philips Imaging DD 001|7a|FL|1|Window Rounding Factor
2001|PHILIPS IMAGING DD 001|7c|US|1|Frame Number
2001|Philips Imaging DD 001|7c|US|1|Frame Number
2001|PHILIPS IMAGING DD 001|80|LO|1|Unknown
2001|Philips Imaging DD 001|80|LO|1|Unknown
2001|PHILIPS IMAGING DD 001|82|IS|1|Echo Train Length
2001|Philips Imaging DD 001|82|IS|1|Echo Train Length
2001|PHILIPS IMAGING DD 001|83|DS|1|Imaging Frequency
2001|Philips Imaging DD 001|83|DS|1|Imaging Frequency
2001|PHILIPS IMAGING DD 001|84|DS|1|Inversion Time
2001|Philips Imaging DD 001|84|DS|1|Inversion Time
2001|PHILIPS IMAGING DD 001|85|DS|1|Magnetic Field Strength
2001|Philips Imaging DD 001|85|DS|1|Magnetic Field Strength
2001|PHILIPS IMAGING DD 001|86|IS|1|Number of Phase Encoding Steps
2001|Philips Imaging DD 001|86|IS|1|Number of Phase Encoding Steps
2001|PHILIPS IMAGING DD 001|87|SH|1|Imaged Nucleus
2001|Philips Imaging DD 001|87|SH|1|Imaged Nucleus
2001|PHILIPS IMAGING DD 001|88|DS|1|Number of Averages
2001|Philips Imaging DD 001|88|DS|1|Number of Averages
2001|PHILIPS IMAGING DD 001|89|DS|1|Phase FOV Percent
2001|Philips Imaging DD 001|89|DS|1|Phase FOV Percent
2001|PHILIPS IMAGING DD 001|8a|DS|1|Sampling Percent
2001|Philips Imaging DD 001|8a|DS|1|Sampling Percent
2001|PHILIPS IMAGING DD 001|8b|SH|1|Transmitting Coil
2001|Philips Imaging DD 001|8b|SH|1|Transmitting Coil
2001|PHILIPS IMAGING DD 001|90|LO|1|Text Foreground Color
2001|Philips Imaging DD 001|90|LO|1|Text Foreground Color
2001|PHILIPS IMAGING DD 001|91|LO|1|Text Background Color
2001|Philips Imaging DD 001|91|LO|1|Text Background Color
2001|PHILIPS IMAGING DD 001|92|LO|1|Text Shadow Color
2001|Philips Imaging DD 001|92|LO|1|Text Shadow Color
2001|PHILIPS IMAGING DD 001|93|LO|1|Text Style
2001|Philips Imaging DD 001|93|LO|1|Text Style
2001|PHILIPS IMAGING DD 001|9a|SQ|1|Unknown
2001|Philips Imaging DD 001|9a|SQ|1|Unknown
2001|PHILIPS IMAGING DD 001|9b|UL|1|Graphic Number
2001|Philips Imaging DD 001|9b|UL|1|Graphic Number
2001|PHILIPS IMAGING DD 001|9c|LO|1|Graphic Annotation Label
2001|Philips Imaging DD 001|9c|LO|1|Graphic Annotation Label
2001|PHILIPS IMAGING DD 001|9f|US|2|Pixel Processing Kernel Size
2001|Philips Imaging DD 001|9f|US|2|Pixel Processing Kernel Size
2001|PHILIPS IMAGING DD 001|a1|CS|1|Is Raw Image
2001|PHILIPS IMAGING DD 001|a3|UL|1|Text Color Foreground
2001|Philips Imaging DD 001|a3|UL|1|Text Color Foreground
2001|PHILIPS IMAGING DD 001|a4|UL|1|Text Color Background
2001|Philips Imaging DD 001|a4|UL|1|Text Color Background
2001|PHILIPS IMAGING DD 001|a5|UL|1|Text Color Shadow
2001|Philips Imaging DD 001|a5|UL|1|Text Color Shadow
2001|PHILIPS IMAGING DD 001|c1|LO|1|Linear Modality GL Transform
2001|Philips Imaging DD 001|c1|LO|1|Linear Modality GL Transform
2001|PHILIPS IMAGING DD 001|c8|LO|1|Exam Card Name
2001|PHILIPS IMAGING DD 001|cc|ST|1|Derivation Description
2001|Philips Imaging DD 001|cc|ST|1|Derivation Description
2001|PHILIPS IMAGING DD 001|da|CS|1|Unknown
2001|Philips Imaging DD 001|da|CS|1|Unknown
2001|PHILIPS IMAGING DD 001|f1|FL|1-n|Prospective Motion Correction
2001|PHILIPS IMAGING DD 001|f2|FL|1-n|Retrospective Motion Correction
2003|Philips X-ray Imaging DD 001|00|CS|1|Unknown
2003|Philips X-ray Imaging DD 001|01|LO|1|Unknown
2003|Philips X-ray Imaging DD 001|02|FD|3|Unknown
2003|Philips X-ray Imaging DD 001|03|LO|1|Unknown
2003|Philips X-ray Imaging DD 001|06|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|09|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|10|LO|1|Unknown
2003|Philips X-ray Imaging DD 001|11|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|12|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|13|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|14|FD|1|Unknown
2003|Philips X-ray Imaging DD 001|15|FD|1|Unknown
2003|Philips X-ray Imaging DD 001|16|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|17|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|18|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|19|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|22|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|24|FD|4|Unknown
2003|Philips X-ray Imaging DD 001|25|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|26|SL|1|Unknown
2003|Philips X-ray Imaging DD 001|27|SH|1|Unknown
2003|Philips X-ray Imaging DD 001|28|SH|1|Unknown
2003|Philips X-ray Imaging DD 001|29|FD|1|Unknown
2003|Philips X-ray Imaging DD 001|2a|LO|1|Unknown
2003|Philips X-ray Imaging DD 001|2b|FD|1|Unknown
2003|Philips X-ray Imaging DD 001|2c|SH|1|Unknown
2003|Philips X-ray Imaging DD 001|2d|SL|1-n|Unknown
2003|Philips X-ray Imaging DD 001|2e|SQ|1|Unknown
2003|Philips X-ray Imaging DD 001|30|CS|1|Unknown
2003|Philips X-ray Imaging DD 001|31|CS|1|Unknown
2003|Philips X-ray Imaging DD 001|32|UI|1|Unknown
2005|PHILIPS MR IMAGING DD 001|00|FL|1|Image Angulation AP
2005|Philips MR Imaging DD 001|00|FL|1|Image Angulation AP
2005|Philips MR Imaging DD 003|00|UL|1|Number of SOP Common
2005|Philips MR Imaging DD 004|00|SS|1|Spectrum Extra Number
2005|Philips MR Imaging DD 005|00|CS|1|Volume View Enabled
2005|PHILIPS MR IMAGING DD 001|01|FL|1|Image Angulation FH
2005|Philips MR Imaging DD 001|01|FL|1|Image Angulation FH
2005|Philips MR Imaging DD 003|01|UL|1|Number of Film Consumption
2005|Philips MR Imaging DD 004|01|SS|1|Spectrum Kx Coordinate
2005|Philips MR Imaging DD 005|01|UL|1|Number of Study Reference
2005|PHILIPS MR IMAGING DD 001|02|FL|1|Image Angulation RL
2005|Philips MR Imaging DD 001|02|FL|1|Image Angulation RL
2005|Philips MR Imaging DD 004|02|SS|1|Spectrum Ky Coordinate
2005|Philips MR Imaging DD 001|03|IS|1|Image Annotation Count
2005|Philips MR Imaging DD 004|03|SS|1|Spectrum Location Number
2005|Philips MR Imaging DD 005|03|UL|1|Number of SPS Codes
2005|PHILIPS MR IMAGING DD 001|04|CS|1|Image Display Orientation
2005|Philips MR Imaging DD 001|04|CS|1|Image Display Orientation
2005|Philips MR Imaging DD 004|04|SS|1|Spectrum Mix Number
2005|Philips MR Imaging DD 005|04|SS|1|Unknown
2005|Philips MR Imaging DD 004|05|SS|1|Spectrum X Coordinate
2005|Philips MR Imaging DD 004|06|SS|1|Spectrum Y Coordinate
2005|Philips MR Imaging DD 005|06|SS|1|Number of PS Specific Character Sets
2005|Philips MR Imaging DD 001|07|IS|1|Image Line Count
2005|Philips MR Imaging DD 004|07|FL|1|Spectrum DC Level
2005|Philips MR Imaging DD 005|07|SS|1|Number of Specific Character Set
2005|PHILIPS MR IMAGING DD 001|08|FL|1|Image Offcenter AP
2005|Philips MR Imaging DD 001|08|FL|1|Image Offcenter AP
2005|Philips MR Imaging DD 004|08|FL|1|Spectrum Noise Level
2005|PHILIPS MR IMAGING DD 001|09|FL|1|Image Offcenter FH
2005|Philips MR Imaging DD 001|09|FL|1|Image Offcenter FH
2005|Philips MR Imaging DD 004|09|FL|1|Spectrum Begin Time
2005|Philips MR Imaging DD 005|09|DS|1|Rescale Intercept Original
2005|PHILIPS MR IMAGING DD 001|0a|FL|1|Image OffCentre RL
2005|Philips MR Imaging DD 001|0a|FL|1|Image OffCentre RL
2005|Philips MR Imaging DD 005|0a|DS|1|Rescale Slope Original
2005|PHILIPS MR IMAGING DD 001|0b|FL|1|Max FP
2005|Philips MR Imaging DD 001|0b|FL|1|Max FP
2005|Philips MR Imaging DD 005|0b|LO|1|Rescale Type Original
2005|PHILIPS MR IMAGING DD 001|0c|FL|1|Min FP
2005|Philips MR Imaging DD 001|0c|FL|1|Min FP
2005|PHILIPS MR IMAGING DD 001|0d|FL|1|Scale Intercept
2005|Philips MR Imaging DD 001|0d|FL|1|Scale Intercept
2005|PHILIPS MR IMAGING DD 001|0e|FL|1|Scale Slope
2005|Philips MR Imaging DD 001|0e|FL|1|Scale Slope
2005|Philips MR Imaging DD 005|0e|SQ|1|Private Shared Sequence
2005|PHILIPS MR IMAGING DD 001|0f|DS|1|Window Center
2005|Philips MR Imaging DD 001|0f|DS|1|Window Center
2005|Philips MR Imaging DD 005|0f|SQ|1|Private Per-Frame Sequence
2005|PHILIPS MR IMAGING DD 001|10|DS|1|Window Width
2005|Philips MR Imaging DD 001|10|DS|1|Window Width
2005|Philips MR Imaging DD 004|10|FL|1|Spectrum Echo Time
2005|Philips MR Imaging DD 005|10|IS|1|MF Conv Treat Spectro Mix Number
2005|PHILIPS MR IMAGING DD 001|11|CS|1|Image Type
2005|Philips MR Imaging DD 001|11|CS|1-n|Image Type
2005|Philips MR Imaging DD 005|11|UI|1|MF Private Referenced SOP Instance UID
2005|PHILIPS MR IMAGING DD 001|12|CS|1|Cardiac Gating
2005|Philips MR Imaging DD 001|12|CS|1|Cardiac Gating
2005|Philips MR Imaging DD 004|12|FL|1|Spectrum Inversion Time
2005|Philips MR Imaging DD 005|12|IS|1|Diffusion B Value Number
2005|PHILIPS MR IMAGING DD 001|13|CS|1|Development Mode
2005|Philips MR Imaging DD 001|13|CS|1|Development Mode
2005|Philips MR Imaging DD 003|13|UL|1|Number of Codes
2005|Philips MR Imaging DD 004|13|SS|1|Spectrum Number
2005|Philips MR Imaging DD 005|13|IS|1|Gradient Orientation Number
2005|PHILIPS MR IMAGING DD 001|14|CS|1|Diffusion
2005|Philips MR Imaging DD 001|14|CS|1|Diffusion
2005|Philips MR Imaging DD 004|14|SS|1|Spectrum Number of Averages
2005|Philips MR Imaging DD 005|14|SL|1|Number of Diffusion B Values
2005|PHILIPS MR IMAGING DD 001|15|CS|1|Fat Saturation
2005|Philips MR Imaging DD 001|15|CS|1|Fat Saturation
2005|Philips MR Imaging DD 002|15|LO|1|User Name
2005|Philips MR Imaging DD 004|15|SS|1|Spectrum Number of Samples
2005|Philips MR Imaging DD 005|15|SL|1|Number of Diffusion Gradient Orientations
2005|PHILIPS MR IMAGING DD 001|16|CS|1|Flow Compensation
2005|Philips MR Imaging DD 001|16|CS|1|Flow Compensation
2005|Philips MR Imaging DD 002|16|LO|1|Pass Word
2005|Philips MR Imaging DD 004|16|SS|1|Spectrum Scan Sequence Number
2005|Philips MR Imaging DD 005|16|CS|1|Plan Mode
2005|PHILIPS MR IMAGING DD 001|17|CS|1|Fourier Interpolation
2005|Philips MR Imaging DD 001|17|CS|1|Fourier Interpolation
2005|Philips MR Imaging DD 002|17|LO|1|Server Name
2005|Philips MR Imaging DD 004|17|SS|1|Spectrum Number of Peaks
2005|Philips MR Imaging DD 005|17|FD|3|Diffusion B Matrix
2005|PHILIPS MR IMAGING DD 001|18|LO|1|Hardcopy Protocol
2005|Philips MR Imaging DD 001|18|LO|1|Hardcopy Protocol
2005|Philips MR Imaging DD 002|18|LO|1|Data Base Name
2005|Philips MR Imaging DD 004|18|SQ|1|Spectrum Peak
2005|Philips MR Imaging DD 005|18|CS|3|Operating Mode Type
2005|PHILIPS MR IMAGING DD 001|19|CS|1|Inverse Reconstructed
2005|Philips MR Imaging DD 001|19|CS|1|Inverse Reconstructed
2005|Philips MR Imaging DD 002|19|LO|1|RootName
2005|Philips MR Imaging DD 004|19|FL|1-n|Spectrum Peak Intensity
2005|Philips MR Imaging DD 005|19|CS|3|Operating Mode
2005|PHILIPS MR IMAGING DD 001|1a|SS|1|Label Syntax
2005|Philips MR Imaging DD 001|1a|SS|1|Label Syntax
2005|Philips MR Imaging DD 005|1a|CS|1|Fat Saturation Technique
2005|PHILIPS MR IMAGING DD 001|1b|CS|1|Magnetization Prepared
2005|Philips MR Imaging DD 001|1b|CS|1|Magnetization Prepared
2005|Philips MR Imaging DD 005|1b|IS|1|Version Number Deleted Images
2005|PHILIPS MR IMAGING DD 001|1c|CS|1|Magnetization Transfer Contrast
2005|Philips MR Imaging DD 001|1c|CS|1|Magnetization Transfer Contrast
2005|Philips MR Imaging DD 005|1c|IS|1|Version Number Deleted Spectra
2005|PHILIPS MR IMAGING DD 001|1d|SS|1|Measurement Scan Resolution
2005|Philips MR Imaging DD 001|1d|SS|1|Measurement Scan Resolution
2005|Philips MR Imaging DD 005|1d|IS|1|Version Number Deleted Blobsets
2005|Philips MR Imaging DD 005|1e|UL|1|LUT1 Offset
2005|Philips MR Imaging DD 005|1f|UL|1|LUT1 Range
2005|Philips MR Imaging DD 002|20|LO|1|DMI Application Name
2005|Philips MR Imaging DD 004|20|LO|1-n|Spectrum Peak Label
2005|Philips MR Imaging DD 005|20|UL|1|LUT1 Begin Color
2005|PHILIPS MR IMAGING DD 001|21|SS|1|Number of Mixes
2005|Philips MR Imaging DD 001|21|SS|1|Number of Mixes
2005|Philips MR Imaging DD 004|21|FL|1-n|Spectrum Peak Phase
2005|Philips MR Imaging DD 005|21|UL|1|LUT1 End Color
2005|PHILIPS MR IMAGING DD 001|22|IS|1|Number of References
2005|Philips MR Imaging DD 001|22|IS|1|Number of References
2005|Philips MR Imaging DD 004|22|FL|1-n|Spectrum Peak Position
2005|Philips MR Imaging DD 005|22|UL|1|LUT2 Offset
2005|PHILIPS MR IMAGING DD 001|23|SS|1|Number of Slabs
2005|Philips MR Imaging DD 001|23|SS|1|Number of Slabs
2005|Philips MR Imaging DD 004|23|CS|1-n|Spectrum Peak Type
2005|Philips MR Imaging DD 005|23|UL|1|LUT2 Range
2005|Philips MR Imaging DD 004|24|FL|1-n|Spectrum Peak Width
2005|Philips MR Imaging DD 005|24|UL|1|LUT2 Begin Color
2005|PHILIPS MR IMAGING DD 001|25|SS|1|Number of Volumes
2005|Philips MR Imaging DD 001|25|SS|1|Number of Volumes
2005|Philips MR Imaging DD 004|25|CS|1|Spectro SI B0 Correction
2005|Philips MR Imaging DD 005|25|UL|1|LUT2 End Color
2005|PHILIPS MR IMAGING DD 001|26|CS|1|Over Sampling Phase
2005|Philips MR Imaging DD 001|26|CS|1|Over Sampling Phase
2005|Philips MR Imaging DD 004|26|FL|1|Spectro B0 Echo Top Position
2005|Philips MR Imaging DD 005|26|CS|1|Viewing Hardcopy Only
2005|PHILIPS MR IMAGING DD 001|27|CS|1|Package Mode
2005|Philips MR Imaging DD 001|27|CS|1|Package Mode
2005|Philips MR Imaging DD 004|27|CS|1|Spectro Complex Component
2005|Philips MR Imaging DD 005|27|CS|1|Unknown
2005|PHILIPS MR IMAGING DD 001|28|CS|1|Partial Fourier Frequency
2005|Philips MR Imaging DD 001|28|CS|1|Partial Fourier Frequency
2005|Philips MR Imaging DD 004|28|CS|1|Spectro Data Origin
2005|Philips MR Imaging DD 005|28|SL|1|Number of Label Types
2005|PHILIPS MR IMAGING DD 001|29|CS|1|PartialFourierPhase
2005|Philips MR Imaging DD 001|29|CS|1|PartialFourierPhase
2005|Philips MR Imaging DD 004|29|FL|1|Spectro Echo Top Position
2005|Philips MR Imaging DD 005|29|CS|1|Label Type
2005|Philips MR Imaging DD 002|2d|LO|1|Root Id
2005|PHILIPS MR IMAGING DD 001|2a|IS|1|Patient Reference ID
2005|Philips MR Imaging DD 001|2a|IS|1|Patient Reference ID
2005|Philips MR Imaging DD 005|2a|CS|1|Exam Print Status
2005|PHILIPS MR IMAGING DD 001|2b|SS|1|Percent Scan Complete
2005|Philips MR Imaging DD 001|2b|SS|1|Percent Scan Complete
2005|Philips MR Imaging DD 005|2b|CS|1|Exam Export Status
2005|PHILIPS MR IMAGING DD 001|2c|CS|1|Phase Encode Reordering
2005|Philips MR Imaging DD 001|2c|CS|1|Phase Encode Reordering
2005|Philips MR Imaging DD 005|2c|CS|1|Exam Storage Commit Status
2005|Philips MR Imaging DD 005|2d|CS|1|Exam Media Write Status
2005|PHILIPS MR IMAGING DD 001|2e|CS|1|PPG PPU Gating
2005|Philips MR Imaging DD 001|2e|CS|1|PPG PPU Gating
2005|Philips MR Imaging DD 005|2e|FL|1|dBdt
2005|PHILIPS MR IMAGING DD 001|2f|CS|1|Spatial Presaturation
2005|Philips MR Imaging DD 001|2f|CS|1|Spatial Presaturation
2005|Philips MR Imaging DD 005|2f|FL|1|Proton SAR
2005|PHILIPS MR IMAGING DD 001|30|FL|1-n|Repetition Time
2005|Philips MR Imaging DD 001|30|FL|1-n|Repetition Time
2005|Philips MR Imaging DD 004|30|CS|1-n|InPlane Transforms
2005|Philips MR Imaging DD 005|30|FL|1|Non Proton SAR
2005|PHILIPS MR IMAGING DD 001|31|CS|1|Respiratory Gating
2005|Philips MR Imaging DD 001|31|CS|1|Respiratory Gating
2005|Philips MR Imaging DD 004|31|SS|1|Number of Spectra Acquired
2005|Philips MR Imaging DD 005|31|FL|1|Local SAR
2005|Philips MR Imaging DD 002|32|SQ|1|Blob Data Object Array
2005|Philips MR Imaging DD 005|32|CS|1|Safety Override Mode
2005|Philips MR Imaging DD 004|33|FL|1|Phase Encoding Echo Top Positions
2005|Philips MR Imaging DD 005|33|DT|1|EV DVD Job In Params Datetime
2005|PHILIPS MR IMAGING DD 001|34|CS|1|Segmented KSpace
2005|Philips MR Imaging DD 001|34|CS|1|Segmented KSpace
2005|Philips MR Imaging DD 002|34|LT|1|Series Transaction UID
2005|Philips MR Imaging DD 003|34|SL|1|Number of Image Per Series Ref
2005|Philips MR Imaging DD 004|34|CS|1|Physical Quantity for Chemical Shift
2005|Philips MR Imaging DD 005|34|DT|1|DVD Job In Params Volume Label
2005|Philips MR Imaging DD 002|35|IS|1|Parent ID
2005|Philips MR Imaging DD 004|35|CS|1|Physical Quantity Spatial
2005|Philips MR Imaging DD 005|35|CS|1|Spectro Examcard
2005|Philips MR Imaging DD 002|36|LO|1|Parent Type
2005|Philips MR Imaging DD 004|36|FL|1|Reference Frequency
2005|Philips MR Imaging DD 005|36|UI|1|Referenced Series Instance UID
2005|PHILIPS MR IMAGING DD 001|37|CS|1|Is Spectro
2005|Philips MR Imaging DD 001|37|CS|1|Is Spectro
2005|Philips MR Imaging DD 002|37|LO|1|Blob Name
2005|Philips MR Imaging DD 004|37|FL|1|Sample Offset
2005|Philips MR Imaging DD 005|37|CS|1|Color LUT Type
2005|PHILIPS MR IMAGING DD 001|38|CS|1|Spoiled
2005|Philips MR Imaging DD 001|38|CS|1|Spoiled
2005|Philips MR Imaging DD 002|38|LO|1|Application Name
2005|Philips MR Imaging DD 004|38|FL|1|Sample Pitch
2005|Philips MR Imaging DD 005|38|LT|1|Unknown
2005|PHILIPS MR IMAGING DD 001|39|CS|1|Steady State
2005|Philips MR Imaging DD 001|39|CS|1|Steady State
2005|Philips MR Imaging DD 002|39|LO|1|Type Name
2005|Philips MR Imaging DD 004|39|SS|2|Search Interval for Peaks
2005|Philips MR Imaging DD 005|39|LT|1|Unknown
2005|PHILIPS MR IMAGING DD 001|3a|SH|1|Sub Anatomy
2005|Philips MR Imaging DD 001|3a|SH|1|Sub Anatomy
2005|Philips MR Imaging DD 005|3a|LT|1|Data Dictionary Contents Version
2005|PHILIPS MR IMAGING DD 001|3b|CS|1|Time Reversed Steady State
2005|Philips MR Imaging DD 001|3b|CS|1|Time Reversed Steady State
2005|Philips MR Imaging DD 005|3b|CS|1|Is Coil Survey
2005|PHILIPS MR IMAGING DD 001|3c|CS|1|Tilt Optimized Nonsaturated Excitation
2005|Philips MR Imaging DD 001|3c|CS|1|Tilt Optimized Nonsaturated Excitation
2005|Philips MR Imaging DD 005|3c|FL|1|Stack Table Position Longitudinal
2005|PHILIPS MR IMAGING DD 001|3d|SS|1|Number of RR Interval Ranges
2005|Philips MR Imaging DD 001|3d|SS|1|Number of RR Interval Ranges
2005|Philips MR Imaging DD 005|3d|FL|1|Stack Table Position Lateral
2005|PHILIPS MR IMAGING DD 001|3e|SL|1-n|RR Intervals Distribution
2005|Philips MR Imaging DD 001|3e|SL|1-n|RR Intervals Distribution
2005|Philips MR Imaging DD 005|3e|FL|1|Stack Posterior Coil Position
2005|PHILIPS MR IMAGING DD 001|3f|SL|1|PlanScan Acquisition Number
2005|Philips MR Imaging DD 001|3f|SL|1|PlanScan Acquisition Number
2005|Philips MR Imaging DD 005|3f|CS|1|Active Implantable Medical Device Limits Applied
2005|Philips MR Imaging DD 001|40|SL|1-n|PlanScan Survey Chemical Shift Number
2005|Philips MR Imaging DD 002|40|LO|1|Version String
2005|Philips MR Imaging DD 004|40|CS|1|Signal Domain for Chemical Shift
2005|Philips MR Imaging DD 005|40|FL|1|Active Implantable Medical Device Head SAR Limit
2005|Philips MR Imaging DD 001|41|SL|1-n|PlanScan Survey Dynamic Scan Number
2005|Philips MR Imaging DD 002|41|LO|1|Comment String
2005|Philips MR Imaging DD 004|41|CS|1|Signal Domain Spatial
2005|Philips MR Imaging DD 005|41|FL|1|Active Implantable Medical Device Whole Body SAR Limit
2005|Philips MR Imaging DD 001|42|SL|1-n|PlanScan Survey Echo Number
2005|Philips MR Imaging DD 002|42|CS|1|Blob In File
2005|Philips MR Imaging DD 004|42|CS|1|Signal Type
2005|Philips MR Imaging DD 005|42|FL|1|Active Implantable Medical Device B1 RMS Limit
2005|Philips MR Imaging DD 001|43|CS|1-n|PlanScan Survey Image Type
2005|Philips MR Imaging DD 002|43|SL|1|Actual Blob Size
2005|Philips MR Imaging DD 003|43|SS|1|No Date of Last Calibration
2005|Philips MR Imaging DD 004|43|CS|1|Spectro Additional Rotations
2005|Philips MR Imaging DD 005|43|FL|1|Active Implantable Medical Device dbDt Limit
2005|Philips MR Imaging DD 001|44|SL|1-n|PlanScan Survey Phase Number
2005|Philips MR Imaging DD 002|44|OW|1|Blob Data
2005|Philips MR Imaging DD 003|44|SS|1|No Time of Last Calibration
2005|Philips MR Imaging DD 004|44|SS|1-n|Spectro Display Ranges
2005|Philips MR Imaging DD 005|44|IS|1|TFE Factor
2005|Philips MR Imaging DD 001|45|SL|1-n|PlanScan Survey Reconstruction Number
2005|Philips MR Imaging DD 002|45|LO|1|Blob Filename
2005|Philips MR Imaging DD 003|45|SS|1|Number of Software Version
2005|Philips MR Imaging DD 004|45|CS|1|Spectro Echo Acquisition
2005|Philips MR Imaging DD 005|45|CS|1|Attenuation Correction
2005|Philips MR Imaging DD 001|46|CS|1-n|PlanScan Survey Scanning Sequence
2005|Philips MR Imaging DD 002|46|SL|1|Blob Offset
2005|Philips MR Imaging DD 004|46|CS|1|Spectro Frequency Unit
2005|Philips MR Imaging DD 005|46|FL|1|FWHM Shim
2005|Philips MR Imaging DD 001|47|SL|1-n|PlanScan Survey Slice Number
2005|Philips MR Imaging DD 002|47|CS|1|Blob Flag
2005|Philips MR Imaging DD 003|47|SS|1|Number of Patient Other Names
2005|Philips MR Imaging DD 004|47|FL|1|Spectro Gamma
2005|Philips MR Imaging DD 005|47|FL|1|Power Optimization
2005|PHILIPS MR IMAGING DD 001|48|IS|1-n|Referenced Acquisition Number
2005|Philips MR Imaging DD 001|48|IS|1-n|Referenced Acquisition Number
2005|Philips MR Imaging DD 003|48|SS|1|Number of Req Recipe of Results
2005|Philips MR Imaging DD 004|48|CS|1|Spectro Hidden Line Removal
2005|Philips MR Imaging DD 005|48|FL|1|Coil Q
2005|PHILIPS MR IMAGING DD 001|49|IS|1-n|Referenced Chemical Shift Number
2005|Philips MR Imaging DD 001|49|IS|1-n|Referenced Chemical Shift Number
2005|Philips MR Imaging DD 003|49|SS|1|Number of Series Operators Name
2005|Philips MR Imaging DD 004|49|FL|1|Spectro Horizontal Shift
2005|Philips MR Imaging DD 005|49|FL|1|Receiver Gain
2005|PHILIPS MR IMAGING DD 001|4a|IS|1-n|Referenced Dynamic Scan Number
2005|Philips MR Imaging DD 001|4a|IS|1-n|Referenced Dynamic Scan Number
2005|Philips MR Imaging DD 005|4a|FL|1|Data Window Duration
2005|PHILIPS MR IMAGING DD 001|4b|IS|1-n|Referenced Echo Number
2005|Philips MR Imaging DD 001|4b|IS|1-n|Referenced Echo Number
2005|Philips MR Imaging DD 005|4b|FL|1|Mixing Time
2005|PHILIPS MR IMAGING DD 001|4c|CS|1-n|Referenced Entity
2005|Philips MR Imaging DD 001|4c|CS|1-n|Referenced Entity
2005|Philips MR Imaging DD 005|4c|FL|1|First Echo Time
2005|PHILIPS MR IMAGING DD 001|4d|CS|1-n|Referenced Image Type
2005|Philips MR Imaging DD 001|4d|CS|1-n|Referenced Image Type
2005|Philips MR Imaging DD 005|4d|CS|1|Is B0 Series
2005|PHILIPS MR IMAGING DD 001|4e|FL|1-n|Slab FOV RL
2005|Philips MR Imaging DD 001|4e|FL|1-n|Slab FOV RL
2005|Philips MR Imaging DD 005|4e|CS|1|Is B1 Series
2005|PHILIPS MR IMAGING DD 001|4f|FL|1-n|Slab Offcentre AP
2005|Philips MR Imaging DD 001|4f|FL|1-n|Slab Offcentre AP
2005|Philips MR Imaging DD 005|4f|CS|1|Volume Select
2005|PHILIPS MR IMAGING DD 001|50|FL|1-n|Slab Offcentre FH
2005|Philips MR Imaging DD 001|50|FL|1-n|Slab Offcentre FH
2005|Philips MR Imaging DD 003|50|SS|1|Number of Series Performing Physicians Name
2005|Philips MR Imaging DD 004|50|FL|2|Spectro Horizontal Window
2005|Philips MR Imaging DD 005|50|SS|1|Number of Patient Other IDs
2005|PHILIPS MR IMAGING DD 001|51|FL|1-n|Slab Offcentre RL
2005|Philips MR Imaging DD 001|51|FL|1-n|Slab Offcentre RL
2005|Philips MR Imaging DD 003|51|SS|1|Number of Study Admitting Diagnostic Description
2005|Philips MR Imaging DD 004|51|SS|1|Spectro Number of Display Ranges
2005|Philips MR Imaging DD 005|51|IS|1|Original Series Number
2005|PHILIPS MR IMAGING DD 001|52|CS|1-n|Slab Type
2005|Philips MR Imaging DD 001|52|CS|1-n|Slab Type
2005|Philips MR Imaging DD 003|52|SS|1|Number of Study Patient Contrast Allergies
2005|Philips MR Imaging DD 004|52|SS|1|Spectro Number of Echo Pulses
2005|Philips MR Imaging DD 005|52|UI|1|Original Series Instance UID
2005|PHILIPS MR IMAGING DD 001|53|CS|1-n|Slab View Axis
2005|Philips MR Imaging DD 001|53|CS|1-n|Slab View Axis
2005|Philips MR Imaging DD 003|53|SS|1|Number of Study Patient Medical Alerts
2005|Philips MR Imaging DD 004|53|LO|1-n|Spectro Processing History
2005|Philips MR Imaging DD 005|53|CS|1|Split Series Job Params
2005|PHILIPS MR IMAGING DD 001|54|FL|1-n|Volume Angulation AP
2005|Philips MR Imaging DD 001|54|FL|1-n|Volume Angulation AP
2005|Philips MR Imaging DD 003|54|SS|1|Number of Study Physicians of Record
2005|Philips MR Imaging DD 004|54|CS|1|Spectro Scan Type
2005|Philips MR Imaging DD 005|54|SS|1|Preferred Dimension for Splitting
2005|PHILIPS MR IMAGING DD 001|55|FL|1-n|Volume Angulation FH
2005|Philips MR Imaging DD 001|55|FL|1-n|Volume Angulation FH
2005|Philips MR Imaging DD 003|55|SS|1|Number of Study Physicians Reading Study
2005|Philips MR Imaging DD 004|55|FL|1-n|Spectro SI CS Intervals
2005|Philips MR Imaging DD 005|55|FD|3|Velocity Encoding Direction
2005|PHILIPS MR IMAGING DD 001|56|FL|1-n|Volume Angulation RL
2005|Philips MR Imaging DD 001|56|FL|1-n|Volume Angulation RL
2005|Philips MR Imaging DD 003|56|SS|1|Number of SC Software Versions
2005|Philips MR Imaging DD 004|56|CS|1|Spectro SI Mode
2005|Philips MR Imaging DD 005|56|SS|1|Contrast/Bolus Number of Injections
2005|PHILIPS MR IMAGING DD 001|57|FL|1-n|Volume FOV AP
2005|Philips MR Imaging DD 001|57|FL|1-n|Volume FOV AP
2005|Philips MR Imaging DD 003|57|SS|1|Number of Running Attributes
2005|Philips MR Imaging DD 004|57|SS|1|Spectro Spectral BW
2005|Philips MR Imaging DD 005|57|LT|1|Contrast/Bolus Agent Code
2005|PHILIPS MR IMAGING DD 001|58|FL|1-n|Volume FOV FH
2005|Philips MR Imaging DD 001|58|FL|1-n|Volume FOV FH
2005|Philips MR Imaging DD 004|58|LO|1|Spectro Title Line
2005|Philips MR Imaging DD 005|58|LT|1|Contrast/Bolus Administration Route Code
2005|PHILIPS MR IMAGING DD 001|59|FL|1-n|Volume FOV RL
2005|Philips MR Imaging DD 001|59|FL|1-n|Volume FOV RL
2005|Philips MR Imaging DD 004|59|FL|1|Spectro Turbo Echo Spacing
2005|Philips MR Imaging DD 005|59|DS|1|Contrast/Bolus Volume
2005|PHILIPS MR IMAGING DD 001|5a|FL|1-n|Volume Offcentre AP
2005|Philips MR Imaging DD 001|5a|FL|1-n|Volume Offcentre AP
2005|Philips MR Imaging DD 005|5a|DS|1|Contrast/Bolus Ingredient Concentration
2005|PHILIPS MR IMAGING DD 001|5b|FL|1-n|Volume Offcentre FH
2005|Philips MR Imaging DD 001|5b|FL|1-n|Volume Offcentre FH
2005|Philips MR Imaging DD 005|5b|IS|1|Contrast/Bolus Dynamic Number
2005|PHILIPS MR IMAGING DD 001|5c|FL|1-n|Volume Offcentre RL
2005|Philips MR Imaging DD 001|5c|FL|1-n|Volume Offcentre RL
2005|Philips MR Imaging DD 005|5c|SQ|1|Contrast/Bolus Sequence
2005|PHILIPS MR IMAGING DD 001|5d|CS|1-n|Volume Type
2005|Philips MR Imaging DD 001|5d|CS|1-n|Volume Type
2005|Philips MR Imaging DD 005|5d|IS|1|Contrast/Bolus ID
2005|PHILIPS MR IMAGING DD 001|5e|CS|1|Volume View Axis
2005|Philips MR Imaging DD 001|5e|CS|1-n|Volume View Axis
2005|PHILIPS MR IMAGING DD 001|60|IS|1|Study Sequence Number
2005|Philips MR Imaging DD 001|60|IS|1|Study Sequence Number
0009|MMCPrivate|1d|SH|1|IsAllowCascadeSave
2005|Philips MR Imaging DD 004|60|FL|1|Spectro Vertical Shift
2005|Philips MR Imaging DD 005|60|CS|1|LUT to RGB Job Params
2005|PHILIPS MR IMAGING DD 001|61|CS|1|Prepulse Type
2005|Philips MR Imaging DD 001|61|CS|1|Prepulse Type
2005|Philips MR Imaging DD 004|61|FL|2|Spectro Vertical Window
2005|Philips MR Imaging DD 004|62|FL|1|Spectro Offset
2005|PHILIPS MR IMAGING DD 001|63|SS|1|fMRI Status Indication
2005|Philips MR Imaging DD 001|63|SS|1|fMRI Status Indication
2005|Philips MR Imaging DD 004|63|FL|1|Spectrum Pitch
2005|PHILIPS MR IMAGING DD 001|64|IS|1-n|Reference Phase Number
2005|Philips MR Imaging DD 001|64|IS|1-n|Reference Phase Number
2005|Philips MR Imaging DD 004|64|CS|1|Volume Selection
2005|PHILIPS MR IMAGING DD 001|65|IS|1-n|Reference Reconstruction Number
2005|Philips MR Imaging DD 001|65|IS|1-n|Reference Reconstruction Number
2005|PHILIPS MR IMAGING DD 001|66|CS|1-n|Reference Scanning Sequence
2005|Philips MR Imaging DD 001|66|CS|1-n|Reference Scanning Sequence
2005|PHILIPS MR IMAGING DD 001|67|IS|1-n|Reference Slice Number
2005|Philips MR Imaging DD 001|67|IS|1-n|Reference Slice Number
2005|PHILIPS MR IMAGING DD 001|68|CS|1-n|Reference Type
2005|Philips MR Imaging DD 001|68|CS|1-n|Reference Type
2005|PHILIPS MR IMAGING DD 001|69|FL|1-n|Slab Angulation AP
2005|Philips MR Imaging DD 001|69|FL|1-n|Slab Angulation AP
2005|PHILIPS MR IMAGING DD 001|6a|FL|1-n|Slab Angulation FH
2005|Philips MR Imaging DD 001|6a|FL|1-n|Slab Angulation FH
2005|PHILIPS MR IMAGING DD 001|6b|FL|1-n|Slab Angulation RL
2005|Philips MR Imaging DD 001|6b|FL|1-n|Slab Angulation RL
2005|PHILIPS MR IMAGING DD 001|6c|FL|1-n|Slab FOV AP
2005|Philips MR Imaging DD 001|6c|FL|1-n|Slab FOV AP
2005|PHILIPS MR IMAGING DD 001|6d|FL|1-n|Slab FOV FH
2005|Philips MR Imaging DD 001|6d|FL|1-n|Slab FOV FH
2005|PHILIPS MR IMAGING DD 001|6e|CS|1-n|Scanning Sequence
2005|Philips MR Imaging DD 001|6e|CS|1-n|Scanning Sequence
2005|PHILIPS MR IMAGING DD 001|6f|CS|1|Acquisition Type
2005|Philips MR Imaging DD 001|6f|CS|1|Acquisition Type
2005|PHILIPS MR IMAGING DD 001|70|LO|1|Hardcopy Protocol EasyVision
2005|Philips MR Imaging DD 001|70|LO|1|Hardcopy Protocol EasyVision
2005|Philips MR Imaging DD 003|70|OW|1|Spectrum Pixel Data
2005|Philips MR Imaging DD 004|70|SS|1|Number Mixes Spectro
2005|PHILIPS MR IMAGING DD 001|71|FL|1-n|Stack Angulation AP
2005|Philips MR Imaging DD 001|71|FL|1-n|Stack Angulation AP
2005|Philips MR Imaging DD 004|71|SQ|1|Series SP Mix
2005|PHILIPS MR IMAGING DD 001|72|FL|1-n|Stack Angulation FH
2005|Philips MR Imaging DD 001|72|FL|1-n|Stack Angulation FH
2005|Philips MR Imaging DD 004|72|SS|40909|SP Mix T Resolution
2005|PHILIPS MR IMAGING DD 001|73|FL|1-n|Stack Angulation RL
2005|Philips MR Imaging DD 001|73|FL|1-n|Stack Angulation RL
2005|Philips MR Imaging DD 004|73|SS|40909|SP Mix KX Resolution
2005|PHILIPS MR IMAGING DD 001|74|FL|1-n|Stack FOV AP
2005|Philips MR Imaging DD 001|74|FL|1-n|Stack FOV AP
2005|Philips MR Imaging DD 004|74|SS|40909|SP Mix KY Resolution
2005|PHILIPS MR IMAGING DD 001|75|FL|1-n|Stack FOV FH
2005|Philips MR Imaging DD 001|75|FL|1-n|Stack FOV FH
2005|Philips MR Imaging DD 004|75|SS|40909|SP Mix F Resolution
2005|PHILIPS MR IMAGING DD 001|76|FL|1-n|Stack FOV RL
2005|Philips MR Imaging DD 001|76|FL|1-n|Stack FOV RL
2005|Philips MR Imaging DD 004|76|SS|40909|SP Mix X Resolution
2005|Philips MR Imaging DD 004|77|SS|40909|SP Mix Y Resolution
2005|PHILIPS MR IMAGING DD 001|78|FL|1-n|Stack Offcentre AP
2005|Philips MR Imaging DD 001|78|FL|1-n|Stack Offcentre AP
2005|Philips MR Imaging DD 004|78|SS|40909|SP Mix Number of Spectra Intended
2005|PHILIPS MR IMAGING DD 001|79|FL|1-n|Stack Offcentre FH
2005|Philips MR Imaging DD 001|79|FL|1-n|Stack Offcentre FH
2005|Philips MR Imaging DD 004|79|SS|40909|SP Mix Number of Averages
2005|PHILIPS MR IMAGING DD 001|7a|FL|1-n|Stack Offcentre RL
2005|Philips MR Imaging DD 001|7a|FL|1-n|Stack Offcentre RL
2005|PHILIPS MR IMAGING DD 001|7b|CS|1-n|Stack Preparation Direction
2005|Philips MR Imaging DD 001|7b|CS|1-n|Stack Preparation Direction
2005|PHILIPS MR IMAGING DD 001|7e|FL|1-n|Stack Slice Distance
2005|Philips MR Imaging DD 001|7e|FL|1-n|Stack Slice Distance
2005|PHILIPS MR IMAGING DD 001|80|SQ|1|Series PlanScan
2005|Philips MR Imaging DD 001|80|SQ|1|Series PlanScan
2005|Philips MR Imaging DD 004|80|SL|1|Number of MF Image Objects
2005|PHILIPS MR IMAGING DD 001|81|CS|1-n|Stack View Axis
2005|Philips MR Imaging DD 001|81|CS|1-n|Stack View Axis
2005|Philips MR Imaging DD 003|81|UI|1|Default Image UID
2005|Philips MR Imaging DD 004|81|IS|1|ScanoGram Survey Number of Images
2005|Philips MR Imaging DD 003|82|CS|1-n|Running Attributes
2005|Philips MR Imaging DD 004|82|UL|1|Number of Procedure Codes
2005|Philips MR Imaging DD 004|83|CS|1-n|Sort Attributes
2005|PHILIPS MR IMAGING DD 001|84|SQ|1|Series Reference
2005|Philips MR Imaging DD 001|84|SQ|1|Series Reference
2005|Philips MR Imaging DD 004|84|SS|1|Number of Sort Attributes
2005|PHILIPS MR IMAGING DD 001|85|SQ|1|Series Volume
2005|Philips MR Imaging DD 001|85|SQ|1|Series Volume
2005|Philips MR Imaging DD 004|85|CS|1|Image Display Direction
2005|PHILIPS MR IMAGING DD 001|86|SS|1|Number of Geometry
2005|Philips MR Imaging DD 001|86|SS|1|Number of Geometry
2005|Philips MR Imaging DD 004|86|CS|1|Inset Scanogram
2005|Philips MR Imaging DD 001|87|SL|1-n|Number of Geometry Slices
2005|Philips MR Imaging DD 004|87|SS|1|Display Layout Number of Columns
2005|Philips MR Imaging DD 001|88|FL|1-n|Geom Angulation AP
2005|Philips MR Imaging DD 004|88|SS|1|Display Layout Number of Rows
2005|Philips MR Imaging DD 001|89|FL|1-n|Geom Angulation FH
2005|Philips MR Imaging DD 004|89|SQ|1|Viewing Protocol
2005|Philips MR Imaging DD 001|8a|FL|1-n|Geom Angulation RL
2005|Philips MR Imaging DD 001|8b|FL|1-n|Geom FOV AP
2005|Philips MR Imaging DD 001|8c|FL|1-n|Geom FOV FH
2005|Philips MR Imaging DD 001|8d|FL|1-n|Geom FOV RL
2005|Philips MR Imaging DD 001|8e|FL|1-n|Geom OffCentre AP
2005|Philips MR Imaging DD 001|8f|FL|1-n|Geom OffCentre FH
2005|Philips MR Imaging DD 001|90|FL|1-n|Geom OffCentre RL
2005|Philips MR Imaging DD 004|90|CS|1|Stack Coil Function
2005|Philips MR Imaging DD 005|90|SQ|1|Original VOI LUT Sequence
2005|Philips MR Imaging DD 001|91|CS|1-n|Geom Preparation Direct
2005|Philips MR Imaging DD 004|91|PN|1|Patient Name Job In Params
2005|Philips MR Imaging DD 005|91|SQ|1|Original Modality LUT Sequence
2005|Philips MR Imaging DD 001|92|FL|1-n|Geom Radial Angle
2005|Philips MR Imaging DD 004|92|IS|1|Geolink ID
2005|Philips MR Imaging DD 001|93|CS|1-n|Geom Radial Axis
2005|Philips MR Imaging DD 004|93|IS|1|Station Number
2005|Philips MR Imaging DD 001|94|FL|1-n|Geom Slice Distance
2005|Philips MR Imaging DD 004|94|CS|1-n|Processing History
2005|Philips MR Imaging DD 001|95|SL|1-n|Geom Slice Number
2005|Philips MR Imaging DD 004|95|UI|1|View Procedure String
2005|Philips MR Imaging DD 001|96|CS|1-n|Geom Type
2005|Philips MR Imaging DD 004|96|CS|1|Flow Images Present
2005|Philips MR Imaging DD 001|97|CS|1-n|Geom ViewA xis
2005|Philips MR Imaging DD 004|97|LO|1|Anatomic Region Code Value
2005|Philips MR Imaging DD 001|98|CS|1-n|Geom Colour
2005|Philips MR Imaging DD 004|98|CS|1|Mobiview Enabled
2005|Philips MR Imaging DD 001|99|CS|1-n|Geom Application Type
2005|Philips MR Imaging DD 002|99|UL|1|Number of Request Excerpts
2005|Philips MR Imaging DD 004|99|CS|1|IViewBold Enabled
2005|Philips MR Imaging DD 001|9a|SL|1-n|Geom Id
2005|Philips MR Imaging DD 001|9b|SH|1-n|Geom Application Name
2005|Philips MR Imaging DD 001|9c|SH|1-n|Geom Label Name
2005|Philips MR Imaging DD 001|9d|CS|1-n|Geom Line Style
2005|PHILIPS MR IMAGING DD 001|9e|SQ|1|Series Geometry
2005|Philips MR Imaging DD 001|9e|SQ|1|Series Geometry
2005|PHILIPS MR IMAGING DD 001|9f|CS|1|Spectral Selective Excitation Pulse
2005|Philips MR Imaging DD 001|9f|CS|1|SeriesSpectral Selective Excitation Pulse
2005|PHILIPS MR IMAGING DD 001|a0|FL|1|Dynamic Scan Begin Time
2005|Philips MR Imaging DD 001|a0|FL|1|Dynamic Scan Begin Time
2005|PHILIPS MR IMAGING DD 001|a2|CS|1|Is COCA
2005|Philips MR Imaging DD 001|a2|CS|1|Is COCA
2005|PHILIPS MR IMAGING DD 001|a3|IS|1|Stack Coil ID
2005|Philips MR Imaging DD 001|a3|IS|1|Stack Coil ID
2005|PHILIPS MR IMAGING DD 001|a4|IS|1|Stack CBB Coil 1
2005|Philips MR Imaging DD 001|a4|IS|1|Stack CBB Coil 1
2005|PHILIPS MR IMAGING DD 001|a5|IS|1|Stack CBB Coil 2
2005|Philips MR Imaging DD 001|a5|IS|1|Stack CBB Coil 2
2005|PHILIPS MR IMAGING DD 001|a6|IS|1|Stack Channel Combination Bitmask
2005|Philips MR Imaging DD 001|a6|IS|1|Stack Channel Combination Bitmask
2005|PHILIPS MR IMAGING DD 001|a7|CS|1|Stack Coil Connection
2005|Philips MR Imaging DD 001|a7|CS|1|Stack Coil Connection
2005|PHILIPS MR IMAGING DD 001|a8|DS|1|Inversion Time
2005|Philips MR Imaging DD 001|a8|DS|1|Inversion Time
2005|PHILIPS MR IMAGING DD 001|a9|CS|1|Geometry Correction
2005|Philips MR Imaging DD 001|a9|CS|1|Geometry Correction
2005|PHILIPS MR IMAGING DD 001|b0|FL|1|Diffusion Direction RL
2005|PHILIPS MR IMAGING DD 001|b1|FL|1|Diffusion Direction AP
2005|PHILIPS MR IMAGING DD 001|b2|FL|1|Diffusion Direction FH
2005|PHILIPS MR IMAGING DD 001|c0|CS|1|Scan Sequence
2005|Philips MR Imaging DD 001|c0|CS|1|Scan Sequence
2007|Philips EV Imaging DD 022|00|ST|1|Unknown
200b|Philips RAD Imaging DD 001|00|PN|1|Unknown
200b|Philips RAD Imaging DD 097|00|ST|1|Unknown
200b|Philips RAD Imaging DD 001|01|US|1|Unknown
200b|Philips RAD Imaging DD 097|01|CS|1|Unknown
200b|Philips RAD Imaging DD 001|02|US|1|Unknown
200b|Philips RAD Imaging DD 097|02|SS|1|Unknown
200b|Philips RAD Imaging DD 001|05|IS|1|Unknown
200b|Philips RAD Imaging DD 001|11|LO|1|Unknown
200b|Philips RAD Imaging DD 001|27|DT|1|Unknown
200b|Philips RAD Imaging DD 001|28|DS|1|Unknown
200b|Philips RAD Imaging DD 001|29|DS|1|Unknown
200b|Philips RAD Imaging DD 001|2a|UL|1|Unknown
200b|Philips RAD Imaging DD 001|2b|DA|1|Unknown
200b|Philips RAD Imaging DD 001|2c|TM|1|Unknown
200b|Philips RAD Imaging DD 001|2d|LO|1|Unknown
200b|Philips RAD Imaging DD 001|3b|LO|1|Unknown
200b|Philips RAD Imaging DD 001|40|SH|1|Unknown
200b|Philips RAD Imaging DD 001|41|SH|1|Unknown
200b|Philips RAD Imaging DD 001|42|UI|1|Unknown
200b|Philips RAD Imaging DD 001|43|UI|1|Unknown
200b|Philips RAD Imaging DD 001|47|DA|1|Unknown
200b|Philips RAD Imaging DD 001|48|SH|1|Unknown
200b|Philips RAD Imaging DD 001|4c|SH|1|Unknown
200b|Philips RAD Imaging DD 001|4d|SH|1|Unknown
200b|Philips RAD Imaging DD 001|4f|DT|1|Unknown
200b|Philips RAD Imaging DD 097|50|SS|1|Unknown
200b|Philips RAD Imaging DD 097|51|SS|1|Unknown
200b|Philips RAD Imaging DD 001|52|CS|1|Unknown
200b|Philips RAD Imaging DD 097|52|SS|1|Unknown
200b|Philips RAD Imaging DD 097|53|SS|1|Unknown
200b|Philips RAD Imaging DD 097|54|ST|1|Unknown
200b|Philips RAD Imaging DD 097|60|LT|1|Unknown
200b|Philips RAD Imaging DD 097|63|LT|1|Unknown
200b|Philips RAD Imaging DD 097|65|SS|1|Unknown
200b|Philips RAD Imaging DD 097|6e|US|1|Unknown
200b|Philips RAD Imaging DD 097|72|FD|1|Unknown
200b|Philips RAD Imaging DD 097|73|SS|1|Unknown
200b|Philips RAD Imaging DD 097|74|IS|1|Unknown
200b|Philips RAD Imaging DD 097|75|CS|1|Unknown
200b|Philips RAD Imaging DD 097|76|SH|1|Unknown
200b|Philips RAD Imaging DD 097|78|IS|1-n|Unknown
200b|Philips RAD Imaging DD 097|79|IS|1|Unknown
200b|Philips RAD Imaging DD 097|7a|IS|1|Unknown
200b|Philips RAD Imaging DD 097|7b|US|1|Unknown
200b|Philips RAD Imaging DD 097|7c|US|1|Unknown
200b|Philips RAD Imaging DD 097|7d|IS|1-n|Unknown
200b|Philips RAD Imaging DD 097|7e|UI|1|Unknown
200b|Philips RAD Imaging DD 097|81|LO|1|Unknown
200b|Philips RAD Imaging DD 097|82|LO|1|Unknown
200b|Philips RAD Imaging DD 097|85|IS|1|Unknown
200b|Philips RAD Imaging DD 097|86|CS|1|Unknown
200b|Philips RAD Imaging DD 097|88|CS|1|Unknown
200b|Philips RAD Imaging DD 097|89|LT|1|Unknown
200b|Philips RAD Imaging DD 097|90|DS|1|Unknown
200b|Philips RAD Imaging DD 097|96|SH|1|Unknown
200b|Philips RAD Imaging DD 097|99|SH|1|Unknown
200b|Philips RAD Imaging DD 097|9a|FD|1|Unknown
200b|Philips RAD Imaging DD 097|9b|FD|1|Unknown
200b|Philips RAD Imaging DD 097|a0|LT|1|Unknown
200d|Philips US Imaging DD 033|00|OB|1|Unknown
200d|Philips US Imaging DD 066|00|OB|1|Unknown
200d|Philips US Imaging DD 109|00|US|1|Unknown
200d|Philips US Imaging DD 033|01|LO|1|Unknown
200d|Philips US Imaging DD 034|01|LO|1|Unknown
200d|Philips US Imaging DD 035|01|LO|1|Unknown
200d|Philips US Imaging DD 038|01|LO|1-n|Unknown
200d|Philips US Imaging DD 039|01|LO|1|Unknown
200d|Philips US Imaging DD 040|01|LO|1|Unknown
200d|Philips US Imaging DD 041|01|LO|1|Unknown
200d|Philips US Imaging DD 048|01|LO|1-n|Unknown
0119|MRSC|1212|IS|1-n|SkeletonizeImage
200d|Philips US Imaging DD 066|01|LO|1|Unknown
200d|Philips US Imaging DD 109|01|SQ|1|Unknown
200d|Philips US Imaging DD 113|01|LO|1|Unknown
200d|Philips US Imaging DD 033|02|LO|1|Unknown
200d|Philips US Imaging DD 034|02|LO|1|Unknown
200d|Philips US Imaging DD 037|02|IS|1|Unknown
200d|Philips US Imaging DD 038|02|LO|1-n|Unknown
200d|Philips US Imaging DD 039|02|LO|1|Unknown
200d|Philips US Imaging DD 040|02|LO|1|Unknown
200d|Philips US Imaging DD 041|02|LO|1|Unknown
200d|Philips US Imaging DD 066|02|LO|1|Unknown
200d|Philips US Imaging DD 109|02|ST|1|Unknown
200d|Philips US Imaging DD 113|02|UL|1|Unknown
200d|Philips US Imaging DD 033|03|LO|1-n|Unknown
200d|Philips US Imaging DD 034|03|LO|1|Unknown
200d|Philips US Imaging DD 035|03|LO|1|Unknown
200d|Philips US Imaging DD 037|03|IS|1|Unknown
200d|Philips US Imaging DD 038|03|LO|1-n|Unknown
200d|Philips US Imaging DD 039|03|LO|1|Unknown
200d|Philips US Imaging DD 040|03|LO|1|Unknown
200d|Philips US Imaging DD 041|03|LO|1|Unknown
200d|Philips US Imaging DD 066|03|LO|1|Unknown
200d|Philips US Imaging DD 109|03|CS|1|Unknown
200d|Philips US Imaging DD 113|03|UL|1|Unknown
200d|Philips US Imaging DD 033|04|LO|1-n|Unknown
200d|Philips US Imaging DD 034|04|LO|1|Unknown
200d|Philips US Imaging DD 035|04|LO|1|Unknown
200d|Philips US Imaging DD 037|04|IS|1|Unknown
200d|Philips US Imaging DD 038|04|LO|1-n|Unknown
200d|Philips US Imaging DD 039|04|LO|1|Unknown
200d|Philips US Imaging DD 040|04|LO|1|Unknown
200d|Philips US Imaging DD 041|04|LO|1|Unknown
200d|Philips US Imaging DD 066|04|LO|1|Unknown
200d|Philips US Imaging DD 109|04|SL|4|Unknown
200d|Philips US Imaging DD 113|04|UL|1|Unknown
200d|Philips US Imaging DD 017|05|LO|1|Unknown
200d|Philips US Imaging DD 033|05|LO|1-n|Unknown
200d|Philips US Imaging DD 034|05|LO|1|Unknown
200d|Philips US Imaging DD 039|05|LO|1|Unknown
200d|Philips US Imaging DD 040|05|LO|1|Unknown
200d|Philips US Imaging DD 043|05|SH|1|Unknown
200d|Philips US Imaging DD 109|05|UL|3|Unknown
200d|Philips US Imaging DD 113|05|UL|1|Unknown
200d|Philips US Imaging DD 033|06|LO|1-n|Unknown
200d|Philips US Imaging DD 037|06|FD|1|Unknown
200d|Philips US Imaging DD 039|06|LO|1|Unknown
200d|Philips US Imaging DD 040|06|LO|1|Unknown
200d|Philips US Imaging DD 041|06|LO|1|Unknown
200d|Philips US Imaging DD 109|06|UL|3|Unknown
200d|Philips US Imaging DD 113|06|UL|1|Unknown
200d|Philips US Imaging DD 021|07|LO|1|Unknown
200d|Philips US Imaging DD 033|07|LO|1|Unknown
200d|Philips US Imaging DD 035|07|LO|1|Unknown
200d|Philips US Imaging DD 039|07|LO|1|Unknown
200d|Philips US Imaging DD 040|07|LO|1|Unknown
200d|Philips US Imaging DD 041|07|LO|1|Unknown
200d|Philips US Imaging DD 065|07|LO|1|Unknown
200d|Philips US Imaging DD 109|07|CS|1|Unknown
200d|Philips US Imaging DD 113|07|CS|1|Unknown
200d|Philips US Imaging DD 033|08|LO|1|Unknown
200d|Philips US Imaging DD 034|08|LO|1|Unknown
200d|Philips US Imaging DD 035|08|LO|1|Unknown
200d|Philips US Imaging DD 037|08|IS|1|Unknown
200d|Philips US Imaging DD 039|08|LO|1|Unknown
200d|Philips US Imaging DD 041|08|LO|1|Unknown
200d|Philips US Imaging DD 109|08|CS|1|Unknown
200d|Philips US Imaging DD 113|08|UL|1|Unknown
200d|Philips US Imaging DD 034|09|LO|1|Unknown
200d|Philips US Imaging DD 035|09|LO|1|Unknown
200d|Philips US Imaging DD 039|09|LO|1|Unknown
200d|Philips US Imaging DD 041|09|LO|1|Unknown
200d|Philips US Imaging DD 043|09|IS|1|Unknown
200d|Philips US Imaging DD 109|09|OB|1|Unknown
200d|Philips US Imaging DD 113|09|UL|1|Unknown
200d|Philips US Imaging DD 034|0a|LO|1|Unknown
200d|Philips US Imaging DD 035|0a|LO|1|Unknown
200d|Philips US Imaging DD 037|0a|IS|1|Unknown
200d|Philips US Imaging DD 039|0a|LO|1|Unknown
200d|Philips US Imaging DD 043|0a|IS|1|Unknown
200d|Philips US Imaging DD 109|0a|UL|1|Unknown
200d|Philips US Imaging DD 113|0a|FD|1|Unknown
200d|Philips US Imaging DD 034|0b|LO|1|Unknown
200d|Philips US Imaging DD 037|0b|LO|1|Unknown
200d|Philips US Imaging DD 039|0b|LO|1|Unknown
200d|Philips US Imaging DD 043|0b|IS|1|Unknown
200d|Philips US Imaging DD 109|0b|OB|1|Unknown
200d|Philips US Imaging DD 113|0b|CS|1|Unknown
200d|Philips US Imaging DD 034|0c|LO|1|Unknown
200d|Philips US Imaging DD 035|0c|LO|1|Unknown
200d|Philips US Imaging DD 037|0c|IS|1|Unknown
200d|Philips US Imaging DD 039|0c|LO|1|Unknown
200d|Philips US Imaging DD 043|0c|IS|1|Unknown
200d|Philips US Imaging DD 109|0c|UL|1|Unknown
200d|Philips US Imaging DD 113|0c|UL|1|Unknown
200d|Philips US Imaging DD 033|0d|LO|1|Private Native Data Type
200d|Philips US Imaging DD 034|0d|LO|1|Unknown
200d|Philips US Imaging DD 035|0d|LO|1|Unknown
200d|Philips US Imaging DD 037|0d|IS|1|Unknown
200d|Philips US Imaging DD 039|0d|LO|1|Unknown
200d|Philips US Imaging DD 043|0d|IS|1|Unknown
200d|Philips US Imaging DD 109|0d|SQ|1|Unknown
200d|Philips US Imaging DD 113|0d|UL|1|Unknown
200d|Philips US Imaging DD 034|0e|LO|1|Unknown
200d|Philips US Imaging DD 037|0e|IS|1|Unknown
200d|Philips US Imaging DD 043|0e|IS|1|Unknown
200d|Philips US Imaging DD 109|0e|CS|1|Unknown
200d|Philips US Imaging DD 113|0e|UL|1|Unknown
200d|Philips US Imaging DD 033|0f|OB|1|Unknown
200d|Philips US Imaging DD 034|0f|LO|1|Unknown
200d|Philips US Imaging DD 037|0f|IS|1|Unknown
200d|Philips US Imaging DD 043|0f|IS|1|Unknown
200d|Philips US Imaging DD 109|0f|LO|1|Unknown
200d|Philips US Imaging DD 113|0f|DS|1|Unknown
200d|Philips US Imaging DD 033|10|IS|1|Private Native Total Num Sample
200d|Philips US Imaging DD 034|10|LO|1|Unknown
200d|Philips US Imaging DD 039|10|LO|1-n|Unknown
200d|Philips US Imaging DD 041|10|LO|1|Unknown
200d|Philips US Imaging DD 043|10|IS|1|Unknown
200d|Philips US Imaging DD 109|10|SL|1|Unknown
200d|Philips US Imaging DD 113|10|DS|1|Unknown
200d|Philips US Imaging DD 033|11|IS|1|Native Data Sample Size
200d|Philips US Imaging DD 034|11|LO|1|Unknown
200d|Philips US Imaging DD 039|11|LO|1-n|Unknown
200d|Philips US Imaging DD 041|11|LO|1|Unknown
200d|Philips US Imaging DD 043|11|IS|1|Unknown
200d|Philips US Imaging DD 109|11|LO|1|Unknown
200d|Philips US Imaging DD 113|11|SL|1|Unknown
200d|Philips US Imaging DD 034|12|LO|1|Unknown
200d|Philips US Imaging DD 039|12|LO|1-n|Unknown
200d|Philips US Imaging DD 041|12|LO|1|Unknown
200d|Philips US Imaging DD 109|12|SL|1|Unknown
200d|Philips US Imaging DD 113|12|UL|1|Unknown
200d|Philips US Imaging DD 034|13|LO|1|Unknown
200d|Philips US Imaging DD 039|13|LO|1-n|Unknown
200d|Philips US Imaging DD 041|13|LO|1|Unknown
200d|Philips US Imaging DD 109|13|US|1-n|Unknown
200d|Philips US Imaging DD 113|13|FL|1-n|Unknown
200d|Philips US Imaging DD 033|14|IS|1|Unknown
200d|Philips US Imaging DD 034|14|LO|1|Unknown
200d|Philips US Imaging DD 039|14|LO|1-n|Unknown
200d|Philips US Imaging DD 041|14|LO|1|Unknown
200d|Philips US Imaging DD 109|14|CS|1|Unknown
200d|Philips US Imaging DD 113|14|SS|1|Unknown
200d|Philips US Imaging DD 033|15|LO|1|Unknown
200d|Philips US Imaging DD 036|15|LO|1-n|Unknown
200d|Philips US Imaging DD 039|15|LO|1|Unknown
200d|Philips US Imaging DD 041|15|LO|1|Unknown
200d|Philips US Imaging DD 042|15|IS|1|Unknown
200d|Philips US Imaging DD 113|15|UL|1|Unknown
200d|Philips US Imaging DD 036|16|LO|1-n|Unknown
200d|Philips US Imaging DD 041|16|LO|1|Unknown
200d|Philips US Imaging DD 042|16|FD|1|Unknown
200d|Philips US Imaging DD 034|17|LO|1|Unknown
200d|Philips US Imaging DD 036|17|LO|1-n|Unknown
200d|Philips US Imaging DD 041|17|LO|1|Unknown
200d|Philips US Imaging DD 043|17|IS|1|Unknown
200d|Philips US Imaging DD 046|17|FD|1|Unknown
200d|Philips US Imaging DD 113|17|FD|1|Unknown
200d|Philips US Imaging DD 034|18|LO|1|Unknown
200d|Philips US Imaging DD 036|18|LO|1-n|Unknown
200d|Philips US Imaging DD 041|18|LO|1|Unknown
200d|Philips US Imaging DD 113|18|FD|1|Unknown
200d|Philips US Imaging DD 036|19|LO|1|Unknown
200d|Philips US Imaging DD 041|19|LO|1|Unknown
200d|Philips US Imaging DD 046|19|LO|1|Unknown
200d|Philips US Imaging DD 113|19|FD|1|Unknown
200d|Philips US Imaging DD 041|1a|LO|1|Unknown
200d|Philips US Imaging DD 043|1a|IS|1|Unknown
200d|Philips US Imaging DD 113|1a|FD|1|Unknown
200d|Philips US Imaging DD 034|1b|LO|1|Unknown
200d|Philips US Imaging DD 041|1b|LO|1|Unknown
200d|Philips US Imaging DD 043|1b|IS|1|Unknown
200d|Philips US Imaging DD 113|1b|FD|1|Unknown
200d|Philips US Imaging DD 034|1c|LO|1|Unknown
200d|Philips US Imaging DD 041|1c|LO|1|Unknown
200d|Philips US Imaging DD 113|1c|FD|1|Unknown
200d|Philips US Imaging DD 034|1d|LO|1|Unknown
200d|Philips US Imaging DD 113|1d|UL|1|Unknown
200d|Philips US Imaging DD 034|1e|LO|1|Unknown
200d|Philips US Imaging DD 043|1e|IS|1|Unknown
200d|Philips US Imaging DD 113|1e|UL|1|Unknown
200d|Philips US Imaging DD 034|1f|LO|1|Unknown
200d|Philips US Imaging DD 043|1f|FD|1|Unknown
200d|Philips US Imaging DD 113|1f|FD|1|Unknown
200d|Philips US Imaging DD 034|20|LO|1|Unknown
200d|Philips US Imaging DD 036|20|LO|1|Unknown
200d|Philips US Imaging DD 040|20|LO|1|Unknown
200d|Philips US Imaging DD 042|20|LO|1|Unknown
200d|Philips US Imaging DD 113|20|FD|1|Unknown
200d|Philips US Imaging DD 033|21|IS|1|Private Native Data Instance Num
200d|Philips US Imaging DD 034|21|LO|1|Unknown
200d|Philips US Imaging DD 043|21|IS|1|Unknown
200d|Philips US Imaging DD 113|21|FD|1|Unknown
200d|Philips US Imaging DD 034|22|LO|1|Unknown
200d|Philips US Imaging DD 113|22|UL|1|Unknown
200d|Philips US Imaging DD 034|23|LO|1|Unknown
200d|Philips US Imaging DD 041|23|LO|1|Unknown
200d|Philips US Imaging DD 043|23|FD|1|Unknown
200d|Philips US Imaging DD 034|24|LO|1|Unknown
200d|Philips US Imaging DD 041|24|LO|1|Unknown
200d|Philips US Imaging DD 043|24|FD|1|Unknown
200d|Philips US Imaging DD 113|24|UL|1|Unknown
200d|Philips US Imaging DD 034|25|LO|1|Unknown
200d|Philips US Imaging DD 041|25|LO|1|Unknown
200d|Philips US Imaging DD 043|25|FD|1|Unknown
200d|Philips US Imaging DD 113|25|UL|1|Unknown
200d|Philips US Imaging DD 034|26|LO|1|Unknown
200d|Philips US Imaging DD 041|26|LO|1|Unknown
200d|Philips US Imaging DD 043|26|FD|1|Unknown
200d|Philips US Imaging DD 113|26|UL|1|Unknown
200d|Philips US Imaging DD 034|27|LO|1|Unknown
200d|Philips US Imaging DD 041|27|LO|1|Unknown
200d|Philips US Imaging DD 043|27|FD|1|Unknown
200d|Philips US Imaging DD 113|27|UL|1|Unknown
200d|Philips US Imaging DD 034|28|LO|1|Unknown
200d|Philips US Imaging DD 041|28|LO|1|Unknown
200d|Philips US Imaging DD 043|28|FD|1|Unknown
200d|Philips US Imaging DD 113|28|UL|1|Unknown
200d|Philips US Imaging DD 041|29|LO|1|Unknown
200d|Philips US Imaging DD 043|29|FD|1|Unknown
200d|Philips US Imaging DD 043|2a|FD|1|Unknown
200d|Philips US Imaging DD 043|2b|FD|1|Unknown
200d|Philips US Imaging DD 043|2c|FD|1-n|Unknown
200d|Philips US Imaging DD 043|2d|FD|1-n|Unknown
200d|Philips US Imaging DD 043|2e|FD|1-n|Unknown
200d|Philips US Imaging DD 043|2f|FD|1-n|Unknown
200d|Philips US Imaging DD 041|30|LO|1|Unknown
200d|Philips US Imaging DD 042|30|LO|1|Unknown
200d|Philips US Imaging DD 043|30|FD|1-n|Unknown
200d|Philips US Imaging DD 042|31|LO|1|Unknown
200d|Philips US Imaging DD 043|31|FD|1-n|Unknown
200d|Philips US Imaging DD 113|31|UL|1|Unknown
200d|Philips US Imaging DD 043|32|FD|1-n|Unknown
200d|Philips US Imaging DD 043|33|FD|1-n|Unknown
200d|Philips US Imaging DD 043|34|FD|1-n|Unknown
200d|Philips US Imaging DD 043|35|IS|1|Unknown
200d|Philips US Imaging DD 043|36|IS|1|Unknown
200d|Philips US Imaging DD 023|37|DA|1|Unknown
200d|Philips US Imaging DD 043|37|FD|1|Unknown
200d|Philips US Imaging DD 023|38|TM|1|Unknown
200d|Philips US Imaging DD 043|38|FD|1-n|Unknown
200d|Philips US Imaging DD 043|39|FD|1|Unknown
200d|Philips US Imaging DD 042|40|LO|1-n|Unknown
200d|Philips US Imaging DD 043|40|IS|1|Unknown
200d|Philips US Imaging DD 043|41|IS|1|Unknown
200d|Philips US Imaging DD 043|42|IS|1|Unknown
200d|Philips US Imaging DD 023|45|IS|1|Unknown
200d|Philips US Imaging DD 039|50|IS|1|Unknown
200d|Philips US Imaging DD 042|50|LO|1-n|Unknown
200d|Philips US Imaging DD 039|51|IS|1|Unknown
200d|Philips US Imaging DD 042|51|LO|1|Unknown
200d|Philips US Imaging DD 039|52|IS|1|Unknown
200d|Philips US Imaging DD 042|52|LO|1|Unknown
200d|Philips US Imaging DD 039|53|IS|1|Unknown
200d|Philips US Imaging DD 042|53|LO|1|Unknown
200d|Philips US Imaging DD 039|54|IS|1|Unknown
200d|Philips US Imaging DD 042|54|LO|1|Unknown
200d|Philips US Imaging DD 039|55|IS|1|Unknown
200d|Philips US Imaging DD 042|55|LO|1|Unknown
200d|Philips US Imaging DD 039|56|IS|1|Unknown
200d|Philips US Imaging DD 042|56|LO|1|Unknown
200d|Philips US Imaging DD 039|57|IS|1|Unknown
200d|Philips US Imaging DD 042|57|LO|1|Unknown
200d|Philips US Imaging DD 039|58|IS|1|Unknown
200d|Philips US Imaging DD 042|58|LO|1|Unknown
200d|Philips US Imaging DD 039|59|IS|1|Unknown
200d|Philips US Imaging DD 042|59|LO|1|Unknown
200d|Philips US Imaging DD 042|5a|LO|1|Unknown
200d|Philips US Imaging DD 042|5b|LO|1|Unknown
200d|Philips US Imaging DD 042|5c|LO|1|Unknown
200d|Philips US Imaging DD 042|5d|LO|1|Unknown
200d|Philips US Imaging DD 042|5e|LO|1|Unknown
200d|Philips US Imaging DD 042|5f|LO|1|Unknown
200d|Philips US Imaging DD 039|60|IS|1|Unknown
200d|Philips US Imaging DD 042|60|LO|1|Unknown
200d|Philips US Imaging DD 039|61|IS|1|Unknown
200d|Philips US Imaging DD 042|70|LO|1|Unknown
200d|Philips US Imaging DD 042|71|LO|1|Unknown
200d|Philips US Imaging DD 042|72|LO|1|Unknown
200d|Philips US Imaging DD 042|73|LO|1|Unknown
200d|Philips US Imaging DD 042|74|LO|1|Unknown
200d|Philips US Imaging DD 042|75|LO|1|Unknown
200d|Philips US Imaging DD 042|76|LO|1|Unknown
200d|Philips US Imaging DD 042|77|LO|1|Unknown
200d|Philips US Imaging DD 042|78|LO|1|Unknown
200d|Philips US Imaging DD 042|8c|LO|1|Unknown
200d|Philips US Imaging DD 045|f1|SQ|1|Unknown
200d|Philips US Imaging DD 045|f3|OB|1|Unknown
200d|Philips US Imaging DD 045|f4|SQ|1|Unknown
200d|Philips US Imaging DD 045|f5|SQ|1|Unknown
200d|Philips US Imaging DD 045|f6|SQ|1|Unknown
200d|Philips US Imaging DD 045|f8|SQ|1|Unknown
200d|Philips US Imaging DD 045|fa|CS|1|Unknown
0009|MMCPrivate|1e|SH|1|IsAllowCascadeProtect
200d|Philips US Imaging DD 045|fb|OB|1|Unknown
4001|Philips Imaging DD 067|00|SQ|1|Unknown
4001|Philips Imaging DD 067|01|CS|1|Unknown
4001|Philips Imaging DD 067|08|CS|1|Unknown
4001|Philips Imaging DD 067|09|CS|1|Unknown
4001|Philips Imaging DD 070|10|SQ|1|Unknown
4001|Philips Imaging DD 070|11|SQ|1|Unknown
4001|Philips Imaging DD 070|12|SQ|1|Unknown
4001|Philips Imaging DD 070|13|ST|1|Unknown
4001|Philips Imaging DD 070|16|ST|1|Unknown
4001|Philips Imaging DD 070|17|ST|1|Unknown
4001|Philips Imaging DD 070|18|ST|1|Unknown
4001|Philips Imaging DD 070|1c|SQ|1|Unknown
4001|Philips Imaging DD 070|1d|LT|1|Unknown
4007|Philips Imaging DD 065|00|CS|1|Unknown
4007|Philips Imaging DD 073|48|FL|1|Unknown
4007|Philips Imaging DD 073|4b|FL|1|Unknown
4007|Philips Imaging DD 073|4c|LO|1|Unknown
4007|Philips Imaging DD 073|4d|FL|1|Unknown
4007|Philips Imaging DD 073|4e|FL|1|Unknown
4007|Philips Imaging DD 073|4f|LO|1|Unknown
7043|Philips NM Private Group|00|SH|1|Unknown
7051|PHILIPS NM -Private|00|US|1|Current Segment
7051|PHILIPS NM -Private|01|US|1|Number of Segments
7051|PHILIPS XCT -Private|01|DS|1|Attenuation Threshold
7051|PHILIPS NM -Private|02|FL|1|Segment Start Position
7051|PHILIPS XCT -Private|02|DS|1|DLPEstimate
7051|PHILIPS NM -Private|03|FL|1|Segment Stop Position
7051|PHILIPS NM -Private|04|FL|1|Relative COR offset - X direction
7051|PHILIPS NM -Private|05|FL|1|Relative COR offset - Z direction
7051|PHILIPS NM -Private|06|US|1|Current Rotation Number
7051|PHILIPS NM -Private|07|US|1|Number of Rotations
7051|PHILIPS NM -Private|10|DS|1-n|Alignment Translations
7051|PHILIPS NM -Private|11|DS|1-n|Alignment Rotations
7051|PHILIPS NM -Private|12|DS|1|Alignment Timestamp
7051|PHILIPS NM -Private|15|UI|1|Related Xray Series Instance UID
7051|PHILIPS NM -Private|25|LO|1|Unknown
7051|PHILIPS NM -Private|26|DS|1|Unknown
7051|PHILIPS NM -Private|27|IS|1|Unknown
7051|PHILIPS NM -Private|28|IS|1|Unknown
7051|PHILIPS NM -Private|29|IS|1|Unknown
7053|Philips PET Private Group|04|OB|1|Unknown
7053|Philips PET Private Group|08|SQ|1|Unknown
7053|Philips PET Private Group|0f|UL|1|Unknown
7053|Philips PET Private Group|10|US|1|Unknown
7053|Philips PET Private Group|11|US|1|Unknown
7053|Philips PET Private Group|12|SQ|1|Unknown
7fe1|SPI-P Release 1|10|OW/OB|1|Pixel Data
7001|Picker NM Private Group|03|OB|1|Unknown
7001|Picker NM Private Group|04|OB|1|Unknown
7001|Picker NM Private Group|05|OB|1|Unknown
7001|Picker NM Private Group|06|OB|1|Unknown
7001|Picker NM Private Group|07|OB|1|Unknown
7001|Picker NM Private Group|08|OB|1|Unknown
7001|Picker NM Private Group|09|OB|1|Unknown
7001|Picker NM Private Group|10|SQ|1|Unknown
7001|Picker NM Private Group|11|LO|1|Unknown
7001|Picker NM Private Group|12|OB|1|Unknown
7001|Picker NM Private Group|13|US|1|Unknown
7001|Picker NM Private Group|14|OB|1|Unknown
7001|Picker NM Private Group|16|OB|1|Unknown
7001|Picker NM Private Group|17|LO|1|Unknown
7101|Picker MR Private Group|00|OB|1|Unknown
7101|Picker MR Private Group|01|SL|1|Unknown
7101|Picker MR Private Group|02|OB|1|Unknown
7101|Picker MR Private Group|03|SL|1|Unknown
7101|Picker MR Private Group|04|SH|1|Unknown
7101|Picker MR Private Group|05|SH|2|Unknown
7101|Picker MR Private Group|06|SH|4|Unknown
7101|Picker MR Private Group|10|DS|1|Unknown
0009|SIEMENS SYNGO INSTANCE MANIFEST|00|SQ|1|Temporary Original Header Sequence
0009|SIEMENS SYNGO INSTANCE MANIFEST|10|AE|1|syngo Index Source AE Title
0009|SIENET|70|DS|1|Unknown
0009|SIENET|71|DS|1|Unknown
0009|SIENET|72|LO|1|Unknown
0009|SIENET|73|LO|1|Unknown
0009|SIENET|74|LO|1|Unknown
0009|SIENET|75|LO|1|Unknown
0009|SIEMENS MED NM|80|ST|1|Unknown
0009|SIEMENS SYNGO INDEX SERVICE|20|DA|1|Object Insertion Date
0009|SIEMENS SYNGO INDEX SERVICE|a0|LO|1|Sender System Device Name
0009|SIEMENS SYNGO INDEX SERVICE|40|DT|1|Last Access Time
0009|SIEMENS SYNGO INDEX SERVICE|41|CS|1|Delete Protected Status
0009|SIEMENS SYNGO INDEX SERVICE|42|CS|1|Received from Archive Status
0009|SIEMENS SYNGO INDEX SERVICE|43|CS|1|Archive Status
0009|SIEMENS SYNGO INDEX SERVICE|44|AE|1|Location
0009|SIEMENS SYNGO INDEX SERVICE|45|CS|1|Logical Deleted Status
0009|SIEMENS SYNGO INDEX SERVICE|46|DT|1|Insert Time
0009|SIEMENS SYNGO INDEX SERVICE|47|IS|1|Visible Instances on Series Level
0009|SIEMENS SYNGO INDEX SERVICE|48|IS|1|Unarchived Instances
0009|SIEMENS SYNGO INDEX SERVICE|49|IS|1|Visible Instances on Study Level
0009|SIEMENS SYNGO INDEX SERVICE|31|SQ|1|Series Object States
0009|SIEMENS SYNGO INDEX SERVICE|30|SQ|1|Instance Object States
0009|SIEMENS SYNGO INDEX SERVICE|50|CS|1|Hidden Instance
0009|SIEMENS AX INSPACE_EP|50|UI|1|Unknown
0009|SIEMENS AX INSPACE_EP|51|UI|1|Unknown
0011|SIEMENS MED NM|10|ST|1|Unknown
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|01|ST|1|Reprocessing Info
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|02|CS|1-n|Data Role Type
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|03|ST|1|Data Role Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|04|SL|1|Rescan Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|05|FD|1|Unknown
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|06|ST|1|Cardiac Type Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|07|ST|1|Cardiac Type Name L2
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|08|ST|1|Misc Indicator
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|09|SL|1|Unknown
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0a|SL|1|Unknown
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0b|DS|1|Unknown
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0c|ST|1|Split Bagging Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0d|ST|1|Split Sub Bagging Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0e|ST|1|Stage Sub Bagging Name
0011|SIEMENS MR DATAMAPPING ATTRIBUTES|0f|ST|1|Is Internal Data Role
0015|ESOFT_DICOM_ECAT_OWNERCODE|00|OB|1|Unknown
0017|SIEMENS MED NM|00|ST|1|Unknown
0017|Siemens: Thorax/Multix FD Version|00|LO|1|Unknown
0017|Siemens: Thorax/Multix FD Version|01|LO|1|Unknown
0017|SIEMENS MED NM|20|ST|1|Unknown
0017|SIEMENS MED NM|70|ST|1|Unknown
0017|SIEMENS MED NM|80|ST|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0a|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0b|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0c|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0d|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0e|LO|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|0f|LO|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|10|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|11|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|14|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|16|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|17|US|1|Unknown
0019|SIEMENS RA PLANE B|b8|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|18|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|19|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|1a|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|1b|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|1c|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|1e|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|1f|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|20|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|21|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|22|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|23|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|24|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|25|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|26|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|27|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|28|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|29|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|48|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|49|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|4d|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|4e|LO|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|4f|LO|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|50|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|51|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|52|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|53|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|54|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|55|SS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|5c|OW|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|64|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|66|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|67|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|68|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|85|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|86|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|87|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|88|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|89|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8a|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8b|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8c|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8d|FL|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8e|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|8f|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a0|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a1|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a2|LO|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a3|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a4|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a5|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|a6|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|aa|US|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|b0|DS|1|Unknown
0017|SIEMENS_FLCOMPACT_VA01A_PROC|c0|LO|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|11|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|12|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|14|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|15|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|16|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|18|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|21|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|22|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|23|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|24|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|25|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|26|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|27|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|2a|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|30|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|31|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|32|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|33|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|37|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|38|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|41|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|43|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|44|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|45|DS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|46|DS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|47|SH|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|48|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|49|LO|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|4a|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|51|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|52|UL|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|61|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|62|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|71|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|72|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|73|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|74|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|79|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|7a|US|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|7b|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|a0|IS|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|c1|LO|1|Unknown
0017|SIEMENS DFR.01 ORIGINAL|c2|LO|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|11|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|12|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|14|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|15|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|25|IS|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|27|IS|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|29|IS|1|Edge Enhancement %
0017|SIEMENS DFR.01 MANIPULATED|30|IS|1|Harmonization %
0017|SIEMENS DFR.01 MANIPULATED|31|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|32|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|33|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|35|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|37|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|38|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|71|IS|1|Landmark
0017|SIEMENS DFR.01 MANIPULATED|72|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|73|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|74|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|77|DS|1|Pixel Shift horizontal
0017|SIEMENS DFR.01 MANIPULATED|78|DS|1|Pixel Shift vertical
0017|SIEMENS DFR.01 MANIPULATED|79|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|7a|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|80|US|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|83|LO|1|Left Marker
0017|SIEMENS DFR.01 MANIPULATED|84|LO|1|Right Marker
0017|SIEMENS DFR.01 MANIPULATED|a1|SH|1|Unknown
0017|SIEMENS DFR.01 MANIPULATED|a2|SH|1|Image Name Extension 1
0017|SIEMENS DFR.01 MANIPULATED|a3|SH|1|Image Name Extension 2
0019|SIEMENS MED SP DXMG WH AWS 1|01|UL|1-n|AEC Coordinates
0019|SIEMENS MED SP DXMG WH AWS 1|02|US|2|AEC Coordinates Size
0019|SIEMENS MED SP DXMG WH AWS 1|10|ST|1|Derivation Description
0019|SIEMENS MED NM|08|SS|1|Unknown
0019|SIEMENS MED NM|0f|SL|1-n|Siemens ICON Data Type
0019|SIEMENS MED NM|16|SS|1|Unknown
0019|SIEMENS MED NM|a5|SS|1-n|Number of Repeats per Phase
0019|SIEMENS MED NM|a6|SS|1-n|Cycles per Repeat
0019|SIEMENS MED NM|a7|SL|1-n|Repeat Start Time
0019|SIEMENS MED NM|a8|SL|1-n|Repeat Stop Time
0019|SIEMENS MED NM|a9|SL|1-n|Effective Repeat Time
0019|SIEMENS MED NM|aa|SS|1-n|Acquired Cycles per Repeat
0019|SIEMENS RA PLANE B|15|OB|1|Unknown
0019|SIEMENS RA PLANE B|ae|UL|1|Unknown
0019|SIEMENS RA PLANE B|b0|US|1|Unknown
0019|SIEMENS RA PLANE B|b1|US|1|Unknown
0019|SIEMENS RA PLANE B|b2|US|1|Unknown
0019|SIEMENS RA PLANE B|b3|US|1|Unknown
0019|SIEMENS RA PLANE B|b4|US|1|Unknown
0019|SIEMENS RA PLANE B|b5|US|1|Unknown
0019|SIEMENS RA PLANE B|b6|US|1|Unknown
0019|SIEMENS RA PLANE B|b7|US|1|Unknown
0019|SIEMENS RA PLANE B|b9|US|1|Unknown
0019|SIEMENS RA PLANE B|bb|UL|1|Unknown
0019|SIEMENS RA PLANE B|bc|UL|1|Unknown
0019|SIEMENS RA PLANE B|bd|UL|1|Unknown
0019|SIEMENS RA PLANE B|be|UL|1|Unknown
0019|SIEMENS RA PLANE B|bf|UL|1|Unknown
0019|SIEMENS RA PLANE B|c0|UL|1|Unknown
0019|SIEMENS RA PLANE B|c1|UL|1|Unknown
0019|SIEMENS RA PLANE B|c2|UL|1|Unknown
0019|SIEMENS RA PLANE B|c3|UL|1|Unknown
0019|SIEMENS RA PLANE B|c4|UL|1|Unknown
0019|SIEMENS RA PLANE B|c5|UL|1|Unknown
0019|SIEMENS RA PLANE B|c6|UL|1|Unknown
0019|SIEMENS RA PLANE B|c7|UL|1|Unknown
0019|SIEMENS RA PLANE B|c8|UL|1|Unknown
0019|SIEMENS RA PLANE B|c9|UL|1|Unknown
0019|SIEMENS RA PLANE B|ca|UL|1|Unknown
0019|SIEMENS RA PLANE B|cb|UL|1|Unknown
0019|SIEMENS RA PLANE B|cc|UL|1|Unknown
0019|SIEMENS RA PLANE B|cd|UL|1|Unknown
0019|SIEMENS RA PLANE B|ce|UL|1|Unknown
0019|SIEMENS RA PLANE B|cf|UL|1|Unknown
0019|SIEMENS RA PLANE B|d1|US|1|Unknown
0019|SIEMENS RA PLANE B|d2|OB|1|Unknown
0019|SIEMENS RA PLANE B|d3|OB|1|Unknown
0019|SIEMENS RA PLANE B|d4|OB|1|Unknown
0019|SIEMENS RA PLANE B|d5|OB|1|Unknown
0019|SIEMENS RA PLANE B|d6|OB|1|Unknown
0019|SIEMENS RA PLANE B|d7|OB|1|Unknown
0019|SIEMENS RA PLANE B|d8|OB|1|Unknown
0019|SIEMENS RA PLANE B|d9|OB|1|Unknown
0019|SIEMENS RA PLANE B|da|OB|1|Unknown
0019|SIEMENS RA PLANE B|db|OB|1|Unknown
0019|SIEMENS RA PLANE B|dc|OB|1|Unknown
0019|SIEMENS RA PLANE B|dd|UL|1|Unknown
0019|SIEMENS RA PLANE B|de|UL|1-n|Unknown
0019|SIEMENS RA PLANE B|df|OB|1|Unknown
0019|SIEMENS RA PLANE B|e0|UL|1|Unknown
0019|SIEMENS CM VA0  CMS|70|DS|1-n|Unknown
0019|SIEMENS CM VA0  CMS|80|LO|1|Unknown
0019|SIEMENS MED NM|93|SL|2|Unknown
0019|SIEMENS CT VA0  COAD|a0|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|a1|DS|1|Unknown
0019|SIEMENS MED NM|a1|SS|1|Unknown
0019|SIEMENS CT VA0  COAD|a2|CS|1|Unknown
0019|SIEMENS CT VA0  COAD|a3|CS|1|Unknown
0019|SIEMENS MED NM|a3|SL|2|Unknown
0019|SIEMENS CT VA0  COAD|a4|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|a5|DS|1|Unknown
0019|SIEMENS CT VA0  COAD|a6|UL|1-n|Unknown
0019|SIEMENS CT VA0  COAD|a7|UL|1-n|Unknown
0019|SIEMENS CT VA0  COAD|a8|UL|1-n|Unknown
0019|SIEMENS CT VA0  COAD|a9|IS|1|Unknown
0019|SIEMENS CT VA0  COAD|aa|CS|1|Unknown
0019|SIEMENS CT VA0  COAD|ab|IS|1|Unknown
0019|SIEMENS CT VA0  COAD|ac|IS|1|Unknown
0019|SIEMENS CT VA0  COAD|ad|IS|1|Unknown
0019|SIEMENS CT VA0  COAD|ae|IS|1|Unknown
0019|SIEMENS CT VA0  COAD|af|DS|1|Unknown
0119|MRSC|1213|IS|1-n|IsotropicResolution
0019|SIEMENS MED NM|c3|ST|1|Unknown
0019|SIEMENS CT VA0  COAD|c4|UL|1|Unknown
0019|SIEMENS CT VA0  COAD|c5|IS|1|Unknown
0019|SIEMENS Selma|06|IS|1|Unknown
0019|SIEMENS Selma|07|IS|1|Unknown
0019|SIEMENS Selma|08|IS|1|Unknown
0019|SIEMENS Selma|26|LO|1|Unknown
0019|SIEMENS Selma|29|LO|1|Unknown
0019|SIEMENS Selma|30|US|1|Unknown
0019|SIEMENS Selma|31|US|1|Unknown
0019|SIEMENS Selma|32|US|1|Unknown
0019|SIEMENS Selma|33|US|1|Unknown
0019|SIEMENS Selma|34|US|1|Unknown
0019|SIEMENS Selma|35|US|1|Unknown
0019|SIEMENS SMS-AX  VIEW 1.0|0a|SS|1|Native Edge Enhancement Kernel Size
0019|SIEMENS SMS-AX  VIEW 1.0|0b|US|1|Subtracted Edge Enhancement Percent Gain
0019|SIEMENS SMS-AX  VIEW 1.0|0c|SS|1|Subtracted Edge Enhancement LUT Index
0019|SIEMENS SMS-AX  VIEW 1.0|0d|SS|1|Subtracted Edge Enhancement Kernel Size
0019|SIEMENS SMS-AX  VIEW 1.0|0e|US|1|Fade Percent
0019|SIEMENS SMS-AX  VIEW 1.0|0f|US|1|Flipped Before Laterality Applied
0019|SIEMENS SMS-AX  VIEW 1.0|11|US|1|Reference Images Taken Flag
0019|SIEMENS SMS-AX  VIEW 1.0|1a|OB|1|Quant 1K Overlay
0019|SIEMENS SMS-AX  VIEW 1.0|1b|US|1|Original Resolution
0019|SIEMENS SMS-AX  VIEW 1.0|1c|DS|1|Auto Window Center
0019|SIEMENS SMS-AX  VIEW 1.0|1d|DS|1|Auto Window Width
0019|SIEMENS SMS-AX  VIEW 1.0|1e|IS|2|Auto Window Correct Value
0019|SIEMENS SMS-AX  VIEW 1.0|1f|DS|1|Sigmoid Window Parameter
0019|SIEMENS SMS-AX  VIEW 1.0|41|SL|2|Dispayed Area Top Left Hand Corner
0019|SIEMENS SMS-AX  VIEW 1.0|42|SL|2|Dispayed Area Bottom Right Hand Corner
0019|SIEMENS SIENET|01|DS|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|00|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|03|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|0c|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|0d|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|0e|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|95|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|20|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|21|FD|1|Unknown
0029|SIEMENS SYNGO VOLUME|44|SQ|1|SubVolume Sequence
0019|SIEMENS CT VA0  COAD|bd|IS|1|Pulmo Trigger Level
0019|SIEMENS CT VA0  COAD|bf|DS|1|Vital Capacity
0019|SIEMENS CT VA0  COAD|c0|DS|1|Pulmo Water
0019|SIEMENS CT VA0  COAD|c1|DS|1|Pulmo Air
0019|SIEMENS CT VA0  COAD|c2|DA|1|Pulmo Date
0019|SIEMENS CT VA0  COAD|c3|TM|1|Pulmo Time
0019|SIEMENS MED SMS USG ANTARES|22|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|23|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|24|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|25|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|26|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|27|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|28|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|29|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|2a|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|2d|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|2e|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|31|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|3a|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|3b|LT|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|40|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|41|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|42|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|43|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|44|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|46|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|47|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|48|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|49|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|54|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|60|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|61|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|62|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|63|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|65|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|66|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|67|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|69|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|6a|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|6c|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|72|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|80|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|81|FD|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|82|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|83|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|86|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|87|SH|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|88|US|1|Unknown
0019|SIEMENS MED SMS USG ANTARES|a0|LT|1|Unknown
0019|Siemens Ultrasound Miscellaneous|20|SH|1|Unknown
0019|Siemens: Thorax/Multix FD Lab Settings|00|LO|1|Unknown
0019|Siemens: Thorax/Multix FD Lab Settings|01|LO|1|Unknown
0029|SIEMENS SYNGO VOLUME|46|UL|1|Histogram Number Of Bins
0019|Siemens: Thorax/Multix FD Lab Settings|02|LO|1|Total Dose Area Product uGy*cm*cm
0019|Siemens: Thorax/Multix FD Lab Settings|03|US|1|Unknown
0019|Siemens: Thorax/Multix FD Lab Settings|04|LO|1|Unknown
0019|Siemens: Thorax/Multix FD Lab Settings|05|US|1|Unknown
0019|Siemens: Thorax/Multix FD Lab Settings|06|FD|1|Table Object Distance
0019|Siemens: Thorax/Multix FD Lab Settings|07|FD|1|Table Detector Distance
0019|Siemens: Thorax/Multix FD Lab Settings|08|US|1-n|Ortho Step Distance
0019|SIEMENS MED SMS USG S2000|00|SH|1|Private Creator Version
0019|SIEMENS MED SMS USG S2000|03|FD|1|Frame Rate
0019|SIEMENS MED SMS USG S2000|0c|US|1|Burned in Graphics
0019|SIEMENS MED SMS USG S2000|0d|SH|1|SieClear Index
0019|SIEMENS MED SMS USG S2000|0e|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|20|SH|1|B-Mode Submode
0019|SIEMENS MED SMS USG S2000|21|FD|1|B-Mode Dynamic Range
0019|SIEMENS MED SMS USG S2000|22|FD|1|B-Mode Overall Gain
0019|SIEMENS MED SMS USG S2000|23|US|1|B-Mode Resolution/Speed Index
0019|SIEMENS MED SMS USG S2000|24|US|1|B-Mode Edge Enhance Index
0019|SIEMENS MED SMS USG S2000|25|US|1|B-Mode Persistence Index
0019|SIEMENS MED SMS USG S2000|26|US|1|B-Mode Map Index
0019|SIEMENS MED SMS USG S2000|27|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|28|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|29|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|2a|US|1|B-Mode Tint Type
0019|SIEMENS MED SMS USG S2000|2d|US|1|B-Mode Tint Index
0019|SIEMENS MED SMS USG S2000|2e|SH|1|ClarifyVE Index
0019|SIEMENS MED SMS USG S2000|30|DS|1|Unknown
0019|SIEMENS MED SMS USG S2000|31|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|3a|US|1|Image Flag
0019|SIEMENS MED SMS USG S2000|3b|LT|1|Unknown
0019|SIEMENS MED SMS USG S2000|40|SH|1|Color Flow State
0019|SIEMENS MED SMS USG S2000|41|US|1|Color Flow Wall Filter Index
0019|SIEMENS MED SMS USG S2000|42|SH|1|Color Flow Submode
0019|SIEMENS MED SMS USG S2000|43|FD|1|Color Flow Overall Gain
0019|SIEMENS MED SMS USG S2000|44|US|1|Color Flow Resolution/Speed Index
0019|SIEMENS MED SMS USG S2000|46|US|1|Color Flow Smooth Index
0019|SIEMENS MED SMS USG S2000|47|US|1|Color Flow Persistence Index
0019|SIEMENS MED SMS USG S2000|48|US|1|Color Flow Map Index
0019|SIEMENS MED SMS USG S2000|49|US|1|Color Flow Priority Index
0019|SIEMENS MED SMS USG S2000|54|FD|1|Color Flow Maximum Velocity
0019|SIEMENS MED SMS USG S2000|60|FD|1|Doppler Dynamic Range
0019|SIEMENS MED SMS USG S2000|61|FD|1|Doppler Overall Gain
0019|SIEMENS MED SMS USG S2000|62|FD|1|Doppler Wall Filter
0019|SIEMENS MED SMS USG S2000|63|FD|1|Doppler Gate Size
0019|SIEMENS MED SMS USG S2000|65|US|1|Doppler Map Index
0029|SIEMENS SYNGO VOLUME|47|OB|1|Volume Histogram Data
0019|SIEMENS MED SMS USG S2000|66|SH|1|Doppler Submode
0019|SIEMENS MED SMS USG S2000|67|US|1|Unknown
0019|SIEMENS MED SMS USG S2000|69|US|1|Doppler Time/Freq Res Index
0019|SIEMENS MED SMS USG S2000|6a|US|1|Doppler Trace Inverted
0019|SIEMENS MED SMS USG S2000|6c|US|1|Doppler Tint Type
0019|SIEMENS MED SMS USG S2000|72|US|1|Doppler Tint Index
0019|SIEMENS MED SMS USG S2000|80|US|1|M-Mode Dynamic Range
0019|SIEMENS MED SMS USG S2000|81|US|1|M-Mode Overall Gain
0019|SIEMENS MED SMS USG S2000|82|US|1|M-Mode Edge Enhance Index
0019|SIEMENS MED SMS USG S2000|83|US|1|M-Mode Map Index
0019|SIEMENS MED SMS USG S2000|86|US|1|M-Mode Tint Type
0019|SIEMENS MED SMS USG S2000|87|SH|1|M-Mode Submode
0019|SIEMENS MED SMS USG S2000|88|US|1|M-Mode Tint Index
0019|SIEMENS MED SMS USG S2000|95|US|1|Unknown
0021|SIEMENS MED NM|00|OB|1|ECAT_Main_Header
0021|SIEMENS MED NM|01|OB|1|ECAT_Image_Subheader
0021|SIEMENS MED ECAT FILE INFO|00|OB|1|ECAT_Main_Header
0021|SIEMENS MED ECAT FILE INFO|01|OB|1|ECAT_Image_Subheader
0021|SIEMENS SMS-AX  ACQ 1.0|09|UL|1|Impac Filename
0021|SIEMENS SMS-AX  ACQ 1.0|0a|UL|1|Copper Filter
0021|SIEMENS SMS-AX  ACQ 1.0|0b|US|1|Measuring Field
0021|SIEMENS SMS-AX  ACQ 1.0|0c|SS|3|Post Blanking Circle
0021|SIEMENS SMS-AX  ACQ 1.0|0d|SS|2-2n|Dyna Angles
0021|SIEMENS SMS-AX  ACQ 1.0|0e|SS|1|Total Steps
0021|SIEMENS SMS-AX  ACQ 1.0|0f|SL|4-n|Dyna X-Ray Info
0021|SIEMENS SMS-AX  ACQ 1.0|1a|US|1|FD Flag
0021|SIEMENS SMS-AX  ACQ 1.0|1b|OB|1|SH_ZOOM
0021|SIEMENS SMS-AX  ACQ 1.0|1c|OB|1|SH_COLPAR
0021|SIEMENS SMS-AX  ACQ 1.0|1d|US|1|K-Factor
0021|SIEMENS SMS-AX  ACQ 1.0|1e|US|8|EVE
0021|SIEMENS SMS-AX  ACQ 1.0|1f|SL|1|Total Scene Time
0021|SIEMENS SMS-AX  ACQ 1.0|27|US|1|IC Stent Flag
0021|SIEMENS SMS-AX  ACQ 1.0|28|SQ|1|Gamma LUT Sequence
0021|SIEMENS SMS-AX  ACQ 1.0|29|DS|1|Acquisition Scene Time
0021|SIEMENS SMS-AX  ACQ 1.0|2a|IS|1|3D Cardiac Phase Center
0021|SIEMENS SMS-AX  ACQ 1.0|2b|IS|1|3D Cardiac Phase Width
0021|SIEMENS SMS-AX  ACQ 1.0|30|OB|1|Organ Program Info
0021|SIEMENS SMS-AX  ACQ 1.0|3a|IS|1|DDO Kernel size
0021|SIEMENS SMS-AX  ACQ 1.0|3b|IS|1|mAs Modulation
0021|SIEMENS SMS-AX  ACQ 1.0|3c|DT|1-n|3D R-Peak Reference Time
0021|SIEMENS SMS-AX  ACQ 1.0|3d|SL|1-n|ECG Frame Time Vector
0021|SIEMENS SMS-AX  ACQ 1.0|3e|SL|1|ECG Start Time of Run
0021|SIEMENS SMS-AX  ACQ 1.0|40|US|3|Gamma LUT Descriptor
0021|SIEMENS SMS-AX  ACQ 1.0|41|LO|1|Gamma LUT Type
0021|SIEMENS SMS-AX  ACQ 1.0|42|US|1-n|Gamma LUT Data
0021|SIEMENS SMS-AX  ACQ 1.0|43|US|1|Global Gain
0021|SIEMENS SMS-AX  ACQ 1.0|44|US|1|Global Offset
0021|SIEMENS SMS-AX  ACQ 1.0|45|US|1|DIPP Mode
0021|SIEMENS SMS-AX  ACQ 1.0|46|US|1|Artis System Type
0021|SIEMENS SMS-AX  ACQ 1.0|47|US|1|Artis Table Type
0021|SIEMENS SMS-AX  ACQ 1.0|48|US|1|Artis Table Top Type
0021|SIEMENS SMS-AX  ACQ 1.0|49|US|1|Water Value
0021|SIEMENS SMS-AX  ACQ 1.0|51|DS|1|3D Positioner Primary Start Angle
0021|SIEMENS SMS-AX  ACQ 1.0|52|DS|1|3D Positioner Secondary Start Angle
0021|SIEMENS SMS-AX  ACQ 1.0|53|SS|3|Stand Position
0021|SIEMENS SMS-AX  ACQ 1.0|54|SS|1|Rotation Angle
0021|SIEMENS SMS-AX  ACQ 1.0|55|US|1|Image Rotation
0021|SIEMENS SMS-AX  ACQ 1.0|56|SS|3|Table Coordinates
0021|SIEMENS SMS-AX  ACQ 1.0|57|SS|3|Isocenter Table Position
0021|SIEMENS SMS-AX  ACQ 1.0|58|DS|1|Table Object Distance
0021|SIEMENS SMS-AX  ACQ 1.0|59|FL|12-n|Carm Coordinate System
0021|SIEMENS SMS-AX  ACQ 1.0|5a|FL|6-n|Robot Axes
0021|SIEMENS SMS-AX  ACQ 1.0|5b|FL|12|Table Coordinate System
0021|SIEMENS SMS-AX  ACQ 1.0|5c|FL|12|Patient Coordinate System
0021|SIEMENS SMS-AX  ACQ 1.0|5d|SS|1-n|Angulation
0021|SIEMENS SMS-AX  ACQ 1.0|5e|SS|1-n|Orbital
0021|SIEMENS SMS-AX  ACQ 1.0|61|SS|1|Large Volume Overlap
0021|SIEMENS SMS-AX  ACQ 1.0|62|US|1|Reconstruction Preset
0021|SIEMENS SMS-AX  ACQ 1.0|63|SS|1|3D Start Angle
0021|SIEMENS SMS-AX  ACQ 1.0|64|SL|1|3D Planned Angle
0021|SIEMENS SMS-AX  ACQ 1.0|65|SL|1|3D Rotation Plane Alpha
0021|SIEMENS SMS-AX  ACQ 1.0|66|SL|1|3D Rotation Plane Beta
0021|SIEMENS SMS-AX  ACQ 1.0|67|SL|1|3D First Image Angle
0021|SIEMENS SMS-AX  ACQ 1.0|68|SS|1-n|3D Trigger Angle
0021|SIEMENS SMS-AX  ACQ 1.0|71|DS|1-n|Detector Rotation
0021|SIEMENS SMS-AX  ACQ 1.0|72|SS|1-n|Physical Detector Rotation
0021|SIEMENS SMS-AX  ACQ 1.0|81|SS|1|Table Tilt
0021|SIEMENS SMS-AX  ACQ 1.0|82|SS|1|Table Rotation
0021|SIEMENS SMS-AX  ACQ 1.0|83|SS|1|Table Cradle Tilt
0021|SIEMENS SMS-AX  ACQ 1.0|a0|OB|1|Crispy1 Container
0021|SIEMENS SMS-AX  ACQ 1.0|a3|SQ|1|3D Cardiac Trigger Sequence
0021|SIEMENS SMS-AX  ACQ 1.0|a4|DT|1|3D Frame Reference Date Time
0021|SIEMENS SMS-AX  ACQ 1.0|a5|FD|1|3D Cardiac Trigger Delay Time
0021|SIEMENS SMS-AX  ACQ 1.0|a6|FD|1|3D R-R Interval Time Measured
0021|Siemens: Thorax/Multix FD Post Processing|00|US|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|01|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|02|FL|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|03|FL|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|04|US|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|05|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|06|FL|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|07|FL|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|08|US|1|Auto Window Flag
0021|Siemens: Thorax/Multix FD Post Processing|09|SL|1|Auto Window Center
0021|Siemens: Thorax/Multix FD Post Processing|0a|SL|1|Auto Window Width
0021|Siemens: Thorax/Multix FD Post Processing|0b|SS|1|Filter ID
0021|Siemens: Thorax/Multix FD Post Processing|0c|FL|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|0d|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|0e|US|1|Dose Control Value
0021|Siemens: Thorax/Multix FD Post Processing|0f|US|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|10|US|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|11|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|12|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|13|SS|1|Unknown
0021|Siemens: Thorax/Multix FD Post Processing|14|US|1|Anatomic Correct View
0021|Siemens: Thorax/Multix FD Post Processing|15|SS|1|Auto Window Shift
0021|Siemens: Thorax/Multix FD Post Processing|16|DS|1|Auto Window Expansion
0021|Siemens: Thorax/Multix FD Post Processing|17|LO|1|System Type
0021|Siemens: Thorax/Multix FD Post Processing|18|LO|1|Detector Type
0021|Siemens: Thorax/Multix FD Post Processing|30|US|1|Anatomic Sort Number
0021|Siemens: Thorax/Multix FD Post Processing|31|US|1|Acquisition Sort Number
0021|SIEMENS MED NM|10|ST|1|Unknown
0021|Siemens: Thorax/Multix FD Lab Settings|08|US|1|Auto Window Flag
0021|Siemens: Thorax/Multix FD Lab Settings|09|SL|1|Auto Window Center
0021|Siemens: Thorax/Multix FD Lab Settings|0a|SL|1|Auto Window Width
0021|Siemens: Thorax/Multix FD Lab Settings|0b|SS|1|Filter ID
0021|Siemens: Thorax/Multix FD Lab Settings|14|US|1|Anatomic Correct View
0021|Siemens: Thorax/Multix FD Lab Settings|15|SS|1|Auto Window Shift
0021|Siemens: Thorax/Multix FD Lab Settings|16|DS|1|Auto Window Expansion
0021|Siemens: Thorax/Multix FD Lab Settings|17|LO|1|System Type
0021|Siemens: Thorax/Multix FD Lab Settings|30|SH|1|Anatomic Sort Number
0021|Siemens: Thorax/Multix FD Lab Settings|31|SH|1|AcquisitionSortNumber
0021|KINETDX_GRAPHICS|a4|OB|1|Unknown
0021|KINETDX|a6|OB|1|Unknown
0021|KINETDX|a5|US|1|Unknown
0021|KINETDX|a8|LO|1|Unknown
0021|KINETDX|aa|OB|1|Unknown
0021|KINETDX|ab|LO|1|Unknown
0021|KINETDX|ac|LO|1|Unknown
0021|KINETDX|b4|LO|1|Unknown
0021|syngoDynamics|ae|OB|1|Unknown
0021|syngoDynamics|b0|LO|1|Unknown
0021|syngoDynamics|b1|LO|1|Unknown
0023|SIEMENS MED NM|01|US|1|DICOM Reader flag
0023|Siemens: Thorax/Multix FD Image Stamp|00|US|1|Unknown
0023|Siemens: Thorax/Multix FD Image Stamp|01|US|1|Unknown
0023|Siemens: Thorax/Multix FD Image Stamp|02|US|1|Unknown
0023|Siemens: Thorax/Multix FD Image Stamp|03|US|1|Unknown
0023|Siemens: Thorax/Multix FD Image Stamp|04|US|1|Unknown
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0a|US|1|Original Number of Frames
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0b|DS|1|Original Scene Duration
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0c|LO|1|Identifier LOID
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0d|SS|1-n|Original Scene VFR Info
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0e|SS|1|Original Frame ECG Position
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|0f|SS|1|Original ECG 1st Frame Offset
0025|SIEMENS SMS-AX  ORIGINAL IMAGE INFO 1.0|16|IS|1|Ready Processing Status
0025|Siemens: Thorax/Multix FD Raw Image Settings|00|SS|1|Raw Image Amplification
0025|Siemens: Thorax/Multix FD Raw Image Settings|01|SS|1|Gamma LUT
0025|Siemens: Thorax/Multix FD Raw Image Settings|02|US|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|03|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|04|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|05|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|06|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|07|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|08|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|09|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|0a|FL|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|0b|US|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|0c|SS|1|Harmonization Kernel
0025|Siemens: Thorax/Multix FD Raw Image Settings|0d|FL|1|Harmonization Gain
0025|Siemens: Thorax/Multix FD Raw Image Settings|0e|SS|1|Edge Enhancement Kernel
0025|Siemens: Thorax/Multix FD Raw Image Settings|0f|FL|1|Edge Enhancement Gain
0025|Siemens: Thorax/Multix FD Raw Image Settings|10|LT|1|Internal Value
0025|Siemens: Thorax/Multix FD Raw Image Settings|11|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|12|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|13|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|14|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|15|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|16|SS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|17|LO|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|18|US|1|Auto Gain
0025|Siemens: Thorax/Multix FD Raw Image Settings|19|US|1|Ortho Subsampling
0009|MMCPrivate|1f|SQ|1|TaskInfo
0025|Siemens: Thorax/Multix FD Raw Image Settings|1a|US|2|Image Crop Upper Left
0025|Siemens: Thorax/Multix FD Raw Image Settings|1b|US|2|Image Crop Upper Right
0025|Siemens: Thorax/Multix FD Raw Image Settings|1c|US|2|Image Crop Lower Left
0025|Siemens: Thorax/Multix FD Raw Image Settings|1d|US|2|Image Crop Lower Right
0025|Siemens: Thorax/Multix FD Raw Image Settings|30|US|1|Manual Cropping
0025|Siemens: Thorax/Multix FD Raw Image Settings|31|SS|1|Gamma LUT Parameter 1
0025|Siemens: Thorax/Multix FD Raw Image Settings|32|DS|1|Gamma LUT Parameter 2
0025|Siemens: Thorax/Multix FD Raw Image Settings|33|SS|1|Gamma LUT Parameter 3
0025|Siemens: Thorax/Multix FD Raw Image Settings|34|SS|1|Gamma LUT Parameter 4
0025|Siemens: Thorax/Multix FD Raw Image Settings|35|LO|1|Gamma LUT Name
0025|Siemens: Thorax/Multix FD Raw Image Settings|36|DS|1|Unknown
0025|Siemens: Thorax/Multix FD Raw Image Settings|37|DS|1|Unknown
0027|SIEMENS SYNGO ENHANCED IDATASET API|01|CS|1|Business Unit Code
0027|SIEMENS SYNGO ENHANCED IDATASET API|02|LO|1|Application Type
0027|SIEMENS SYNGO ENHANCED IDATASET API|03|SQ|1|Application Attributes Sequence
0029|SIEMENS SYNGO FUNCTION ASSIGNMENT|01|LO|1|Data Reference
0029|SHS MagicView 300|02|FD|1|Unknown
0029|SHS MagicView 300|03|FD|1|Unknown
0029|SIEMENS MED DISPLAY|80|US|1|Unknown
0029|SIEMENS MED MAMMO|5a|CS|1|Unknown
0029|SIEMENS MED DISPLAY 0000|99|CS|1|Unknown
0029|SIEMENS MED DISPLAY 0000|c1|US|1-n|Unknown
0029|SIEMENS MED DISPLAY 0000|b0|US|1|Unknown
0029|SIEMENS MED DISPLAY 0000|b2|US|1-n|Unknown
0029|SIEMENS MED DISPLAY 0001|99|CS|1|Unknown
0029|SIEMENS MED DISPLAY 0001|a0|US|1|Unknown
0029|SIEMENS MED DISPLAY 0001|a1|US|1|Unknown
0029|SIEMENS MED DISPLAY 0001|a2|US|1-n|Unknown
0119|MRSC|1220|IS|1-n|MedianFilterKernel
0029|SIEMENS MEDCOM HEADER|77|UL|1|Referenced Object Offset
0029|SIEMENS SYNGO VOLUME|12|US|1|Slices
0029|SIEMENS SYNGO VOLUME|14|OB|1|Volume Histogram
0029|SIEMENS SYNGO VOLUME|18|IS|1|Volume Level
0029|SIEMENS SYNGO VOLUME|30|DS|3|Voxel Spacing
0029|SIEMENS SYNGO VOLUME|32|DS|3|Volume Position (Patient)
0029|SIEMENS SYNGO VOLUME|37|DS|9|Volume Orientation (Patient)
0029|SIEMENS SYNGO VOLUME|40|CS|1|Resampling Flag
0029|SIEMENS SYNGO VOLUME|42|CS|1|Normalization Flag
0029|SIEMENS MEDCOM HEADER|71|AT|1|Referenced Tag
0029|SIEMENS MEDCOM HEADER|72|CS|1|Referenced Tag Type
0029|SIEMENS MEDCOM HEADER|73|UL|1|Referenced Value Length
0029|SIEMENS MEDCOM HEADER|74|CS|1|Referenced Object Device Type
0029|SIEMENS MEDCOM HEADER|76|OB|1|Referenced Object ID
0029|SIEMENS SYNGO TIME POINT SERVICE|01|LO|1|Time Point ID
0029|SIEMENS SYNGO TIME POINT SERVICE|02|LO|1|Time Point Information
0029|SIEMENS SYNGO TIME POINT SERVICE|50|SQ|1|Studies in Time Point Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|00|CS|1|Presentation Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|01|CS|1|Presentation Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|02|SQ|1|Advanced Presentation Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|03|SQ|1|Time Point Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|04|SQ|1|Base Image Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|05|SQ|1|Overlay Image Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|06|SQ|1|Registration Instance Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|07|SQ|1|Real World Value Mapping Instance Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|08|SQ|1|Measurement Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|09|UI|1|Measurement UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|10|SQ|1|Segmentation Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|11|UI|1|Segmentation UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|12|SQ|1|Navigation Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|13|CS|1|Navigation Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|14|CS|1|Auto Navigation Direction
0029|SIEMENS SYNGO ADVANCED PRESENTATION|15|DS|1|Auto Navigation Frame Rate
0029|SIEMENS SYNGO ADVANCED PRESENTATION|16|CS|1|Auto Navigation Mode
0029|SIEMENS SYNGO ADVANCED PRESENTATION|17|DS|1|Auto Navigation Realtime Speed
0029|SIEMENS SYNGO ADVANCED PRESENTATION|18|CS|1|Auto Navigation Strategy
0029|SIEMENS SYNGO ADVANCED PRESENTATION|19|CS|1|Auto Navigation Realtime Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|20|IS|1|Index Navigation Current Index
0029|SIEMENS SYNGO ADVANCED PRESENTATION|21|IS|1|Index Auto Navigation Skipping Degree
0029|SIEMENS SYNGO ADVANCED PRESENTATION|22|DS|1|Volume Navigation Minimum Pixel Spacing
0029|SIEMENS SYNGO ADVANCED PRESENTATION|23|CS|1|Volume Navigation Scroll Unit
0029|SIEMENS SYNGO ADVANCED PRESENTATION|24|DS|1|Volume Navigation Step Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|25|DS|1|Volume Navigation Jump Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|26|IS|1|Referenced Registration Number
0029|SIEMENS SYNGO ADVANCED PRESENTATION|27|UI|1|Real World Value Mapping UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|28|DS|1|Channel Alpha Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|30|LO|1|Measurement Application Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|31|SQ|1|Measurement Data Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|32|LO|1|Measurement Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|33|UI|1|Measurement Frame of Reference UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|34|UI|1|Measurement UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|35|IS|1|Measurement Application Number
0029|SIEMENS SYNGO ADVANCED PRESENTATION|36|ST|1|Measurement Application Number Prefix Text
0029|SIEMENS SYNGO ADVANCED PRESENTATION|37|CS|1|Measurement Graphic Is Visible Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|38|UI|4|Referenced Syngo UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|39|UI|1|Clinical Finding UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3a|CS|1|Measurement Evaluation String Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3b|IS|1|Measurement Evaluation Integer Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3c|FL|1|Measurement Evaluation Decimal Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3d|CS|1|Measurement Line Show Center Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3e|CS|1|Measurement Angle Show ArrowTip Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|3f|SQ|1|Camera Home Settings Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|40|DS|1|Camera Zoom
0029|SIEMENS SYNGO ADVANCED PRESENTATION|41|DS|3|Camera Position
0029|SIEMENS SYNGO ADVANCED PRESENTATION|42|DS|4|Camera Orientation
0029|SIEMENS SYNGO ADVANCED PRESENTATION|43|DS|1|Camera Far Clip Plane
0029|SIEMENS SYNGO ADVANCED PRESENTATION|44|DS|1|Camera Near Clip Plane
0029|SIEMENS SYNGO ADVANCED PRESENTATION|45|DS|1|Camera Thickness
0029|SIEMENS SYNGO ADVANCED PRESENTATION|46|DS|1|Camera ViewPort Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|47|DS|1|Camera Aspect Ratio
0029|SIEMENS SYNGO ADVANCED PRESENTATION|48|LO|1|Camera Projection Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|49|DS|1|Camera Field of View
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4a|DS|1|Camera Image Plane Distance
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4b|DS|1|Camera Image Maximum Height
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4c|DS|1|Camera Image Minimum Height
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4d|DS|1|Parallel Shift Interval MM
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4e|DS|3|Parallel Shift BoundingBox Minimum
0029|SIEMENS SYNGO ADVANCED PRESENTATION|4f|DS|3|Parallel Shift BoundingBox Maximum
0029|SIEMENS SYNGO ADVANCED PRESENTATION|50|CS|1|Renderer Vertex Is Characteristic Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|51|CS|1|Renderer Thickness Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|52|DS|4|Renderer Threshold
0029|SIEMENS SYNGO ADVANCED PRESENTATION|53|DS|4|Renderer Material
0029|SIEMENS SYNGO ADVANCED PRESENTATION|54|DS|4|Renderer DirectionalLight Color
0029|SIEMENS SYNGO ADVANCED PRESENTATION|55|DS|3|Renderer DirectionalLight Direction
0029|SIEMENS SYNGO ADVANCED PRESENTATION|56|CS|1|Renderer DirectionalLight TwoSide Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|57|SQ|1|Renderer PWL TransferFunction Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|58|IS|0-n|Renderer PWL Vertex Index
0029|SIEMENS SYNGO ADVANCED PRESENTATION|59|DS|0-n|Renderer PWL Vertex Color
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5a|CS|1|Renderer Is Camera Required Flag
0119|MRSC|1221|DS|1-n|BackgroundCorrection
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5b|CS|1|Renderer Do Depth Test Flag 
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5c|CS|1|Renderer Directional Light Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5d|SQ|1|Renderer Thickness Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5e|SQ|0-n|Renderer Slice Spacing Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|5f|DS|1|Renderer Sampling Distance
0029|SIEMENS SYNGO ADVANCED PRESENTATION|60|DS|1|Renderer Initial Sampling Distance
0029|SIEMENS SYNGO ADVANCED PRESENTATION|61|SQ|1|Segmentation Display Data Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|62|UI|0-n|Segmentation Display Data UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|63|SQ|1|Segmentation Display Parameter Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|64|LO|1|Segmentation Display Parameter Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|65|LO|1|Segmentation Display Visibility
0029|SIEMENS SYNGO ADVANCED PRESENTATION|66|DS|4|Segmentation Display Color
0029|SIEMENS SYNGO ADVANCED PRESENTATION|67|CS|1|Segmentation Display is Selected Flag 
0029|SIEMENS SYNGO ADVANCED PRESENTATION|68|OB|1|Segmentation Additional Information Blob
0029|SIEMENS SYNGO ADVANCED PRESENTATION|69|ST|1|Hash Code Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|6a|LO|1-n|Segmentation Version Identifier
0029|SIEMENS SYNGO ADVANCED PRESENTATION|70|DS|3|Segmentation Volume Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|71|UI|1-n|Registration Referenced Frames
0029|SIEMENS SYNGO ADVANCED PRESENTATION|72|UI|1-n|Registration Referenced Registrations
0029|SIEMENS SYNGO ADVANCED PRESENTATION|73|LO|1|Registration Creation Algorithm Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|74|CS|1|ECG Graphic Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|7a|DS|1|Segmentation Volume Storage Data Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|7b|FL|16|Segmentation Volume Model Matrix
0029|SIEMENS SYNGO ADVANCED PRESENTATION|80|DS|3|Camera Rotation Axis
0029|SIEMENS SYNGO ADVANCED PRESENTATION|81|SL|0-n|Overlay Hidden Display Attributes
0029|SIEMENS SYNGO ADVANCED PRESENTATION|82|LO|1|Presentation State Group Identifier
0029|SIEMENS SYNGO ADVANCED PRESENTATION|83|US|1|Temporary Smallest Image Pixel Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|84|DS|3|Camera Rotation Center
0029|SIEMENS SYNGO ADVANCED PRESENTATION|85|CS|1|Camera Rotation Center Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|86|DS|12|Camera Parallel Epiped
0029|SIEMENS SYNGO ADVANCED PRESENTATION|87|DS|1|Camera Max Zoom In Factor
0029|SIEMENS SYNGO ADVANCED PRESENTATION|88|DS|1|Camera Min Zoom In Factor
0029|SIEMENS SYNGO ADVANCED PRESENTATION|89|US|1|Temporary Largest Image Pixel Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|8a|CS|1|Camera Rotation Axis Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|8b|DS|3|Measurement Surface Normal
0029|SIEMENS SYNGO ADVANCED PRESENTATION|8c|FL|16|Measurement Ellipsoid Model Matrix
0029|SIEMENS SYNGO ADVANCED PRESENTATION|8d|LO|1|Measurement Evaluation DataRole ID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|8e|LO|1|Measurement Algorithm Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|91|SQ|1|Measurement Evaluation DataRole Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|92|CS|1|Measurement Evaluation DataRole Item
0029|SIEMENS SYNGO ADVANCED PRESENTATION|93|SQ|1|Measurement Evaluation Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|94|DS|1|Measurement Evaluation Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|95|CS|1|Measurement Evaluation ID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|96|FL|0-n|Measurement Data Points
0029|SIEMENS SYNGO ADVANCED PRESENTATION|97|FL|0-n|Measurement Data Angles
0029|SIEMENS SYNGO ADVANCED PRESENTATION|98|LO|1|Measurement Data Slice
0029|SIEMENS SYNGO ADVANCED PRESENTATION|99|FL|1|Measurement Data Slice Thickness
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9a|SQ|1|Measurement Referenced Frames Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9b|DS|0-n|Measurement Evaluation Longest Distance
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9c|DS|0-n|Measurement Evaluation Centroid
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9d|FL|6|Measurement Data Bounding Box 
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9e|LO|1|Measurement Text
0029|SIEMENS SYNGO ADVANCED PRESENTATION|9f|IS|1|Measurement Diameter
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a0|DS|1|Image Rotation Fractional
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a1|LO|1|Preset Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a2|SQ|1|Fusion LUT Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a3|CS|1|Fusion LUT Is Active Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a5|UI|1|Syngo UID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a6|UI|1|Presentation Version Identifier
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a7|SQ|1|Presentation Module Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a8|LO|1|Presentation Module Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|a9|SQ|1|Presentation State Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|aa|CS|1|LUT Inverted Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ab|IS|1|Softcopy VOI LUT Viewing Index
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ac|FD|2|Displayed Area Bottom Right Hand Corner Fractional
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ad|FD|2|Displayed Area Top Left Hand Corner Fractional
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ae|FL|1|Measurement Alpha
0029|SIEMENS SYNGO ADVANCED PRESENTATION|af|OB|1|Measurement Bitmap
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b0|US|1|Current Frame Number
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b1|LO|1|Image Text View Name
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b2|SQ|1|Image Text View Content Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b3|LO|1-n|Image Text Line Names
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b4|LO|1-n|ImageText Line Values
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b5|SQ|1|Measurement Evaluation Text Position Sequence
0033|SIEMENS MED NM|1a|FL|1-n|Unknown
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b6|CS|1|Measurement Link Evaluation Text Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b7|DS|3|Measurement Evaluation Text Position Vector
0029|SIEMENS SYNGO ADVANCED PRESENTATION|b8|OB|1|Image Text Alpha Blending Line Value
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c1|SQ|1|Task Data Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c2|CS|1|Task Data Type
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c3|LO|1|Task Data Version
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c4|ST|1|Task Data Description
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c5|OB|1|Task Data
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c6|IS|1|Task Data Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|c9|SQ|1|Clip Plane Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ca|DS|3|Clip Plane Center
0029|SIEMENS SYNGO ADVANCED PRESENTATION|cb|DS|3|Clip Plane Normal
0029|SIEMENS SYNGO ADVANCED PRESENTATION|cc|DS|2|Clip Plane Scale
0029|SIEMENS SYNGO ADVANCED PRESENTATION|cd|CS|1|Clip Plane Use Thickness Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|ce|DS|1|Clip Plane Thickness
0029|SIEMENS SYNGO ADVANCED PRESENTATION|cf|SQ|1|Image Sequence
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d0|CS|1|Clip Plane Enable Clip
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d1|DS|1|Clip Plane Handle Ratio
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d2|DS|24|Clip Plane Bounding Points
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d3|DS|16|Clip Plane Motion Matrix
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d4|DS|1|Clip Plane Shift Velocity
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d5|CS|1|Clip Plane Enabled Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d6|DS|1|Clip Plane Rotate Velocity
0029|SIEMENS SYNGO ADVANCED PRESENTATION|d7|CS|1|Clip Plane Show Graphics Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|e0|DS|3|Crop Box Size
0029|SIEMENS SYNGO ADVANCED PRESENTATION|e1|CS|1|Crop Box Enabled Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|e2|DS|3|Crop Box Absolute Origin
0029|SIEMENS SYNGO ADVANCED PRESENTATION|e3|CS|1|Crop Box Show Graphics Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f1|DS|0-n|Curved Camera Coordinates
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f2|DS|1|Curved Camera Point of Interest
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f3|CS|1|Curved Camera Point of Interest Usage Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f4|DS|1|Curved Camera Thickness
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f5|DS|1|Curved Camera Extrusion Length
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f6|CS|1|Curved Camera Rotation Axis Mode
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f7|DS|1|Curved Camera Roll Rotation Axis
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f8|DS|1|Curved Camera View Port Height
0029|SIEMENS SYNGO ADVANCED PRESENTATION|f9|DS|1|Curved Camera Cut Direction
0029|SIEMENS SYNGO ADVANCED PRESENTATION|fa|DS|1|Curved Camera Pan Vector
0029|SIEMENS SYNGO ADVANCED PRESENTATION|fb|LO|1|Clinical Finding ID
0029|SIEMENS SYNGO ADVANCED PRESENTATION|fc|CS|1|Measurement Is Circle Flag
0029|SIEMENS SYNGO ADVANCED PRESENTATION|fd|LO|1|Measurement Application Type ID
0029|SIEMENS SYNGO FRAME SET|10|SQ|1|Image Frame Sequence
0029|SIEMENS SYNGO FRAME SET|12|CS|1|Type of Progression
0029|SIEMENS SYNGO FRAME SET|14|IS|1|Representation Level
0029|SIEMENS SYNGO FRAME SET|16|SQ|1|Representation Information Sequence
0029|SIEMENS SYNGO FRAME SET|18|IS|1|Number of Representations
0029|SIEMENS SYNGO FRAME SET|20|IS|1|Representation Pixel Offset
0029|SIEMENS SYNGO PRINT SERVICE|10|IS|1|Sheet Number
0029|SIEMENS IKM CKS LUNGCAD BMK|01|UT|1|Unknown
0029|SIEMENS IKM CKS CXRCAD FINDINGS|01|UT|1|Unknown
0029|SIEMENS MED NM|08|CS|1|Modality Image Header Type
0029|SIEMENS MED NM|09|LO|1|Modality Image Header Version
0029|SIEMENS MED NM|10|OB|1|Modality Image Header Info
0031|SIEMENS MED NM|01|ST|1|Unknown
0031|SIEMENS MED NM|0c|SS|1|Unknown
0031|SIEMENS MED NM|0f|SL|1|Unknown
0031|SIEMENS MED NM|10|SL|1|Unknown
0031|SIEMENS MED NM|12|SS|1|Unknown
0031|SIEMENS MED NM|13|ST|1|Unknown
0031|SIEMENS MED NM|14|ST|1|Unknown
0031|SIEMENS MED NM|15|SL|1-n|Unknown
0031|SIEMENS MED NM|16|SL|1-n|Unknown
0031|SIEMENS MED NM|17|SS|1-n|Unknown
0031|SIEMENS MED NM|20|ST|1|Unknown
0031|SIEMENS MED NM|21|SS|1|Unknown
0031|SIEMENS SYNGO SOP CLASS PACKING|10|SQ|1|SOP Class Packing Sequence
0031|SIEMENS SYNGO SOP CLASS PACKING|20|CS|1|Packing Version
0031|SIEMENS SYNGO SOP CLASS PACKING|21|CS|1|Packing Originator
0031|SIEMENS SYNGO SOP CLASS PACKING|30|UI|1|Original SOP Class UID
0031|SIEMENS SYNGO SOP CLASS PACKING|31|UI|1|Original Study Instance UID
0031|SIEMENS SYNGO SOP CLASS PACKING|32|UI|1|Original Series Instance UID
0031|SIEMENS SYNGO SOP CLASS PACKING|33|UI|1|Original SOP Instance UID
0031|SIEMENS SYNGO SOP CLASS PACKING|34|UI|1|Original Transfer Syntax UID
0031|SIEMENS SYNGO SOP CLASS PACKING|40|AT|1-n|Attributes to Set to Zero Length
0031|SIEMENS SYNGO SOP CLASS PACKING|41|AT|1-n|Attributes to Remove
0031|SIEMENS SYNGO SOP CLASS PACKING|50|US|1|Original Rows
0031|SIEMENS SYNGO SOP CLASS PACKING|51|US|1|Original Columns
0031|SIEMENS SYNGO SOP CLASS PACKING|58|CS|2-n|Original Image Type
0031|SIEMENS SYNGO SOP CLASS PACKING|60|CS|1|Original Modality
0029|SIEMENS CSA ENVELOPE|11|OB|1|syngo Report Presentation
0029|SIEMENS CSA REPORT|08|CS|1|Report Type
0029|SIEMENS CSA REPORT|09|LO|1|Report Version
0029|SIEMENS CSA REPORT|15|US|1|SR Variant
0029|SIEMENS CSA REPORT|17|UI|1|SC SOP Instance UID
0033|SIEMENS MED NM|20|FL|1|Bed correction angle
0031|SIEMENS SYNGO SOP CLASS PACKING|70|SQ|1|Sequence of Original StreamCchunks
0031|SIEMENS SYNGO SOP CLASS PACKING|71|AT|1|Start Tag of a Stream Chunk
0031|SIEMENS SYNGO SOP CLASS PACKING|72|AT|1|End Tag of a Stream Chunk
0031|SIEMENS SYNGO SOP CLASS PACKING|73|CS|1|Stream Chunk is a Payload
0031|SIEMENS SYNGO SOP CLASS PACKING|80|OB|1|Stream Chunk
0031|SIEMENS SYNGO WORKFLOW|10|UI|1|Internal Patient UID
0031|SIEMENS SYNGO WORKFLOW|11|SH|1|Patients Death Indicator
0031|SIEMENS SYNGO WORKFLOW|12|DA|1|Patients Death Date
0031|SIEMENS SYNGO WORKFLOW|13|TM|1|Patients Death Time
0031|SIEMENS SYNGO WORKFLOW|14|SH|1|VIP Indicator
0031|SIEMENS SYNGO WORKFLOW|15|US|1|Emergency Flag
0031|SIEMENS SYNGO WORKFLOW|20|SH|1|Internal Visit UID
0031|SIEMENS SYNGO WORKFLOW|25|SH|1|Internal ISR UID
0031|SIEMENS SYNGO WORKFLOW|32|SH|1|Control State
0031|SIEMENS SYNGO WORKFLOW|34|US|1|Local Flag
0031|SIEMENS SYNGO WORKFLOW|36|UI|1-n|Referenced Studies
0031|SIEMENS SYNGO WORKFLOW|40|LO|1|Workflow ID
0031|SIEMENS SYNGO WORKFLOW|41|LO|1|Workflow Description
0031|SIEMENS SYNGO WORKFLOW|42|LO|1|Workflow Control State
0031|SIEMENS SYNGO WORKFLOW|43|US|1|Workflow Ad Hoc Flag
0031|SIEMENS SYNGO WORKFLOW|44|US|1|Hybrid Flag
0031|SIEMENS SYNGO WORKFLOW|50|LO|1|Workitem ID
0031|SIEMENS SYNGO WORKFLOW|51|LO|1|Workitem Name
0031|SIEMENS SYNGO WORKFLOW|52|LO|1|Workitem Type
0031|SIEMENS SYNGO WORKFLOW|53|LO|1-n|Workitem Roles
0031|SIEMENS SYNGO WORKFLOW|54|LO|1|Workitem Description
0031|SIEMENS SYNGO WORKFLOW|55|LO|1|Workitem Control State
0031|SIEMENS SYNGO WORKFLOW|56|LO|1|Claiming User
0031|SIEMENS SYNGO WORKFLOW|57|LO|1|Claiming Host
0031|SIEMENS SYNGO WORKFLOW|58|LO|1|Taskflow ID
0031|SIEMENS SYNGO WORKFLOW|59|LO|1|Taskflow Name
0031|SIEMENS SYNGO WORKFLOW|5a|US|1|Failed Flag
0031|SIEMENS SYNGO WORKFLOW|5b|DT|1|Scheduled Time
0031|SIEMENS SYNGO WORKFLOW|5c|US|1|Workitem Ad Hoc Flag
0031|SIEMENS SYNGO WORKFLOW|5d|US|1|Patient Update Pending Flag
0031|SIEMENS SYNGO WORKFLOW|5e|US|1|Patient Mixup Flag
0031|SIEMENS SYNGO WORKFLOW|60|LO|1|Client ID
0031|SIEMENS SYNGO WORKFLOW|61|LO|1|Template ID
0031|SIEMENS SYNGO WORKFLOW|81|LO|1|Institution Name
0031|SIEMENS SYNGO WORKFLOW|82|ST|1|Institution Address
0031|SIEMENS SYNGO WORKFLOW|83|SQ|1|Institution Code Sequence
0119|MRSC|1222|DS|1-n|UnSharpMasking
0033|SIEMENS MED NM|01|FL|1-n|Flood Correction Matrix Detector 2
0033|SIEMENS MED NM|10|FL|1-n|COR Data for Detector 1
0033|SIEMENS MED NM|11|FL|1-n|COR Data for Detector 2
0033|SIEMENS MED NM|14|FL|1|MHR ( Y-Shift) data for detector 1
0033|SIEMENS MED NM|15|FL|1|MHR ( Y-Shift) data for detector 2
0033|SIEMENS MED NM|18|FL|1-n|NCO Data for detector 1
0119|MRSC|1223|IS|1-n|LocalThresholdKernel
0037|SIEMENS MED NM|00|OW|1|Flood correction matrix Detector 1
0037|SIEMENS MED NM|80|OW|1|Flood correction matrix Detector 2
0041|SIEMENS MED SP DXMG WH AWS 1|02|SH|1|Reason for the Requested Procedure
0041|SIEMENS MED NM|30|ST|1|Unknown
0041|SIEMENS MED NM|32|ST|1|Unknown
0041|SIEMENS MI RWVM SUV|01|CS|1|SUV Decay Correction Method
0051|SIEMENS MED SP DXMG WH AWS 1|10|DS|1|Unknown
0051|SIEMENS MED SP DXMG WH AWS 1|37|DS|6|Unknown
0051|SIEMENS MED SP DXMG WH AWS 1|50|UI|1|Unknown
0033|SIEMENS MED NM|22|SS|1-n|Bed U/D correction data
0033|SIEMENS MED NM|23|SS|1-n|Gantry L/R Correction Data
0033|SIEMENS MED NM|24|FL|1|BackProjection Correction angle head 1
0033|SIEMENS MED NM|25|FL|1|BackProjection Correction angle head 2
0033|SIEMENS MED NM|28|SL|1|MHR calibrations
0033|SIEMENS MED NM|29|FL|1-n|Crystal thickness
0033|SIEMENS MED NM|30|LO|1|Preset name used for acquisition
0033|SIEMENS MED NM|31|FL|1|Camera Config Angle
0033|SIEMENS MED NM|32|LO|1|Crystal Type
0033|SIEMENS MED NM|33|SL|1|Coin Gantry Step
0033|SIEMENS MED NM|34|FL|1|Wholebody bed step
0033|SIEMENS MED NM|36|FL|1|Coincidence weight factor table
0033|SIEMENS MED NM|37|SL|1|Starburst flags at image acq time
0033|SIEMENS MED NM|38|FL|1|Pixel Scale factor
0035|SIEMENS MED NM|00|LO|1|Specialized Tomo Type
0035|SIEMENS MED NM|01|LO|1|Energy Window Type
0035|SIEMENS MED NM|02|SS|1|Start and End Row Illuminated By Wind Position
0035|SIEMENS MED NM|03|LO|1|Blank Scan Image For Profile
0035|SIEMENS MED NM|04|SS|1|Repeat Number of the Original Dynamic SPECT
0035|SIEMENS MED NM|05|SS|1|Phase Number of the Original Dynamic SPECT
0035|SIEMENS MED NM|06|LO|1|Siemens Profile 2 Image Subtype
0039|SIEMENS MED NM|00|LT|1|Toshiba CBF Activity Results
0039|SIEMENS MED NM|01|LT|1|Related CT Series Instance UID
0041|SIEMENS MED NM|01|SL|1|Whole Body Tomo Position Index
0041|SIEMENS MED NM|02|SL|1|Whole Body Tomo Number of Positions
0041|SIEMENS MED NM|03|FL|1|Horizontal Table Position of CT scan
0041|SIEMENS MED NM|04|FL|1|Effective Energy fo CT Scan
0041|SIEMENS MED NM|05|FD|1-n|Long Linear Drive Information for Detector 1
0041|SIEMENS MED NM|06|FD|1-n|Long Linear Drive Information for Detector 2
0041|SIEMENS MED NM|07|FD|1-n|Trunnion Information for Detector 1
0041|SIEMENS MED NM|08|FD|1-n|Trunnion Information for Detector 2
0041|SIEMENS MED NM|09|FL|1|Broad Beam Factor
0041|SIEMENS MED NM|0a|FD|1|Original Wholebody Position
0041|SIEMENS MED NM|0b|FD|1|Wholebody Scan Range
0041|SIEMENS MED NM|10|FL|40910|Effective Emission Energy
0041|SIEMENS MED NM|11|FL|1-n|Gated Frame Duration
0043|SIEMENS MED NM|01|FL|1-n|Detector View Angle
0043|SIEMENS MED NM|02|FD|40923|Transformation Matrix
0043|SIEMENS MED NM|04|FL|1-n|View Dependent Y Shift MHR For Detector 2
0045|SIEMENS MED NM|01|LO|1-n|Planar Processing String
0051|SIEMENS MED SP DXMG WH AWS 1|60|DS|1|Primary Positioner Scan Arc
0051|SIEMENS MED SP DXMG WH AWS 1|61|DS|1|Secondary Positioner Scan Arc
0051|SIEMENS MED SP DXMG WH AWS 1|62|DS|1|Primary Positioner Scan Start Angle
0051|SIEMENS MED SP DXMG WH AWS 1|63|DS|1|Secondary Positioner Scan Start Angle
0051|SIEMENS MED SP DXMG WH AWS 1|64|DS|1|Primary Positioner Increment
0051|SIEMENS MED SP DXMG WH AWS 1|65|DS|1|Secondary Positioner Increment
0055|SIEMENS MED NM|20|SS|1|Unknown
0055|SIEMENS MED NM|22|SS|1|Unknown
0055|SIEMENS MED NM|24|SS|1|Unknown
0055|SIEMENS MED NM|30|SS|1|Unknown
0055|SIEMENS MED NM|32|SS|1|Unknown
0055|SIEMENS MED NM|34|SS|1|Unknown
0055|SIEMENS MED NM|40|SS|1|Unknown
0055|SIEMENS MED NM|42|SS|1|Unknown
0055|SIEMENS MED NM|44|SS|1|Unknown
0055|SIEMENS MED NM|4c|SL|1|Unknown
0055|SIEMENS MED NM|4d|SL|1|Unknown
0055|SIEMENS MED NM|51|SS|1|Unknown
0055|SIEMENS MED NM|52|SS|1|Unknown
0055|SIEMENS MED NM|53|ST|1|Unknown
0055|SIEMENS MED NM|55|SL|1|Unknown
0055|SIEMENS MED NM|5c|ST|1|Unknown
0055|SIEMENS MED NM|6d|SS|1|Unknown
0055|SIEMENS MED NM|a8|SS|1|Unknown
0055|SIEMENS MED NM|c2|SS|1|Unknown
0055|SIEMENS MED NM|c3|SS|1|Unknown
0055|SIEMENS MED NM|c4|SS|1|Unknown
0055|SIEMENS MED NM|d0|SS|1|Unknown
0055|SIEMENS MED SP DXMG WH AWS 1|01|LO|1|Projection View Display String
0055|SIEMENS MED NM|05|SS|1|Random Window Width
0055|SIEMENS MED NM|7e|FL|2|Collimator Thickness mm
0055|SIEMENS MED NM|7f|FL|2|Collimator Angular Resolution radians
0055|SIEMENS MED NM|c0|SS|1-n|Useful Field of View
0057|SIEMENS MED NM|02|FL|1|Dose Calibration Factor
0057|SIEMENS MED NM|03|LO|1|Units
0057|SIEMENS MED NM|04|LO|1|Decay Correction
0057|SIEMENS MED NM|05|SL|1-n|Radionuclide Half Life
0057|SIEMENS MED NM|06|FL|1|Rescale Intercept
0057|SIEMENS MED NM|07|FL|1|Rescale Slope
0057|SIEMENS MED NM|08|FL|1|Frame Reference Time
0057|SIEMENS MED NM|09|SL|1|Number of Radiopharmaceutical Information Sequence
0057|SIEMENS MED NM|0a|FL|1|Decay Factor
0057|SIEMENS MED NM|0b|LO|1|Counts Source
0057|SIEMENS MED NM|0c|SL|1-n|Radionuclide Positron Fraction
0057|SIEMENS MED NM|0e|US|1-n|Trigger Time of CT Slice
0061|SIEMENS MED NM|01|FL|1-n|X Principal Ray Offset
0061|SIEMENS MED NM|05|FL|1-n|Y Principal Ray Offset
0061|SIEMENS MED NM|09|FL|1-n|X Principal Ray Angle
0061|SIEMENS MED NM|0a|FL|1-n|Y Principal Ray Angle
0061|SIEMENS MED NM|0b|FL|1-n|X Short Focal Length
0061|SIEMENS MED NM|0c|FL|1-n|Y Short Focal Length
0061|SIEMENS MED NM|0d|FL|1-n|X Long Focal Length
0061|SIEMENS MED NM|0e|FL|1-n|Y Long Focal Length
0119|MRSC|1224|IS|1-n|AbsoluteLimits
0071|SIEMENS WH SR 1.0|01|LO|1|Unknown
0071|SIEMENS WH SR 1.0|02|LO|1|Unknown
0071|SIEMENS MED PT|23|US|1|Volume Index
0071|SIEMENS MED PT|24|IS|1|Time Slice Duration
0071|SIEMENS SYNGO REGISTRATION|20|SQ|1|Registered Image Sequence
0071|SIEMENS SYNGO REGISTRATION|21|CS|1|Registration Is Validated Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|00|SQ|1|Graphic Object Sequence
0061|SIEMENS MED NM|10|FL|1-n|Y Focal Scaling
0061|SIEMENS MED NM|11|FL|1-n|X Motion Correction Shift
0061|SIEMENS MED NM|15|FL|1-n|Y Motion Correction Shift
0061|SIEMENS MED NM|19|FL|1|X Heart Center
0061|SIEMENS MED NM|1a|FL|1|Y Heart Center
0061|SIEMENS MED NM|1b|FL|1|Z Heart Center
0061|SIEMENS MED NM|1c|LO|1|Image Pixel Content Type
0061|SIEMENS MED NM|1d|SS|1|Auto Save Corrected Series
0061|SIEMENS MED NM|1e|LT|1|Distorted Series Instance UID
0061|SIEMENS MED NM|21|SS|1-n|Recon Range
0061|SIEMENS MED NM|22|LO|1|Recon Orientation
0061|SIEMENS MED NM|24|FL|1|Recon Transverse Angle
0061|SIEMENS MED NM|25|FL|1|Recon Sagittal Angle
0061|SIEMENS MED NM|26|FL|1|Recon X Mask Size
0061|SIEMENS MED NM|27|FL|1|Recon Y Mask Size
0061|SIEMENS MED NM|28|FL|1|Recon X Image Center
0061|SIEMENS MED NM|29|FL|1|Recon Y Image Center
0061|SIEMENS MED NM|2a|FL|1|Recon Z Image Center
0061|SIEMENS MED NM|2b|FL|1|Recon X Zoom
0061|SIEMENS MED NM|2c|FL|1|Recon Y Zoom
0061|SIEMENS MED NM|2d|FL|1|Recon Threshold
0061|SIEMENS MED NM|2e|FL|1|Recon Output Pixel Size
0061|SIEMENS MED NM|2f|LO|1-n|Scatter Estimation Method
0061|SIEMENS MED NM|30|LO|1-n|Scatter Estimation Method Mode
0061|SIEMENS MED NM|31|FL|1-n|Scatter Estimation Lower Window Weights
0061|SIEMENS MED NM|32|FL|1-n|Scatter Estimation Upper Window Weights
0061|SIEMENS MED NM|33|LO|1-n|Scatter Estimation Window Mode
0061|SIEMENS MED NM|34|LO|1-n|Scatter Estimation Filter
0061|SIEMENS MED NM|35|LO|1|Recon RawTomo Input UID
0061|SIEMENS MED NM|36|LO|1|Recon CT Input UID
0061|SIEMENS MED NM|37|FL|1|Recon Z Mask Size
0061|SIEMENS MED NM|38|FL|1|Recon X Mask Center
0061|SIEMENS MED NM|39|FL|1|Recon Y Mask Center
0061|SIEMENS MED NM|3a|FL|1|Recon Z Mask Center
0061|SIEMENS MED NM|51|LT|1|Raw Tomo Series UID
0061|SIEMENS MED NM|53|LT|1|HighRes CT Series UID
0071|SIEMENS MED PT WAVEFORM|46|UN|1|Starting Respiratory Amplitude
0071|SIEMENS MED PT WAVEFORM|47|UN|1|Starting Respiratory Phase
0071|SIEMENS MED PT WAVEFORM|48|UN|1|Ending Respiratory Amplitude
0071|SIEMENS MED PT WAVEFORM|49|UN|1|Ending Respiratory Phase
0071|SIEMENS MED PT WAVEFORM|50|CS|1|Respiratory Trigger Type
0071|SIEMENS MED PT|21|UI|1|Registration Matrix UID
0071|SIEMENS MED PT|22|DT|1|Decay Correction DateTime
0071|SIEMENS SYNGO OBJECT GRAPHICS|01|SL|1|Fill Style Version
0071|SIEMENS SYNGO OBJECT GRAPHICS|02|FL|4|Fill Background Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|03|FL|4|Fill Foreground Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|04|SL|1|Fill Mode
0071|SIEMENS SYNGO OBJECT GRAPHICS|05|OB|1|Fill Pattern
0071|SIEMENS SYNGO OBJECT GRAPHICS|06|SL|1|Line Style Version
0071|SIEMENS SYNGO OBJECT GRAPHICS|07|FL|4|Line Background Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|08|FL|4|Line Foreground Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|09|DS|1|Line Type
0071|SIEMENS SYNGO OBJECT GRAPHICS|10|DS|1|Line Thickness
0071|SIEMENS SYNGO OBJECT GRAPHICS|11|DS|1|Line Shadow X Offset
0071|SIEMENS SYNGO OBJECT GRAPHICS|12|DS|1|Line Shadow Y Offset
0071|SIEMENS SYNGO OBJECT GRAPHICS|13|DS|1|Shadow Style
0071|SIEMENS SYNGO OBJECT GRAPHICS|14|FL|4|Shadow Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|15|DS|1|Stipple Pattern
0071|SIEMENS SYNGO OBJECT GRAPHICS|16|DS|1|Line Anti Aliasing
0071|SIEMENS SYNGO OBJECT GRAPHICS|17|CS|1|Line-Z-Blend Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|18|SL|1|Text Style Version
0071|SIEMENS SYNGO OBJECT GRAPHICS|19|FL|4|Text Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|20|SL|1|Text Horizontal Align
0071|SIEMENS SYNGO OBJECT GRAPHICS|21|SL|1|Text Vertical Align
0071|SIEMENS SYNGO OBJECT GRAPHICS|22|DS|1|Text Shadow X Offset
0071|SIEMENS SYNGO OBJECT GRAPHICS|23|DS|1|Text Shadow Y Offset
0071|SIEMENS SYNGO OBJECT GRAPHICS|24|SL|1|Text Shadow Style
0071|SIEMENS SYNGO OBJECT GRAPHICS|25|FL|4|Text Shadow Color
0071|SIEMENS SYNGO OBJECT GRAPHICS|26|CS|1-n|Text Log Font
0071|SIEMENS SYNGO OBJECT GRAPHICS|27|CS|1|Text-Z-Blend Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|28|OB|1|Graphic Bit Mask
0071|SIEMENS SYNGO OBJECT GRAPHICS|29|CS|1|Visiblility Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|30|SL|1|Graphic Sensitivity
0071|SIEMENS SYNGO OBJECT GRAPHICS|31|SL|1|Graphic Pick Mode Type
0071|SIEMENS SYNGO OBJECT GRAPHICS|32|SL|1|Graphic Layer
0071|SIEMENS SYNGO OBJECT GRAPHICS|33|SL|1|Graphic Object Version
0071|SIEMENS SYNGO OBJECT GRAPHICS|34|SL|1|Graphic Coordinate System
0071|SIEMENS SYNGO OBJECT GRAPHICS|35|CS|1|Graphic Custom Attributes
0071|SIEMENS SYNGO OBJECT GRAPHICS|36|CS|1|Graphic Custom Attributes Key
0071|SIEMENS SYNGO OBJECT GRAPHICS|37|CS|1|Graphic Custom Attributes Value
0071|SIEMENS SYNGO OBJECT GRAPHICS|38|CS|1|Graphic View Name
0071|SIEMENS SYNGO OBJECT GRAPHICS|39|DS|3|Graphic Data
0071|SIEMENS SYNGO OBJECT GRAPHICS|40|CS|1|Graphic Type
0071|SIEMENS SYNGO OBJECT GRAPHICS|41|US|1|Number of Graphic Points
0071|SIEMENS SYNGO OBJECT GRAPHICS|42|DS|1|Axis Main Tick Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|43|DS|1|Axis Detail Tick Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|44|DS|1|Axis Main Tick Spacing
0071|SIEMENS SYNGO OBJECT GRAPHICS|45|DS|1-n|Axis Detail Tick Spacing
0071|SIEMENS SYNGO OBJECT GRAPHICS|46|DS|1|Axis Main Tick Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|47|DS|1|Axis Detail Tick Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|48|SL|1|Axis Tick Behavior
0071|SIEMENS SYNGO OBJECT GRAPHICS|49|SL|1|Axis Tick Aligment
0071|SIEMENS SYNGO OBJECT GRAPHICS|50|DS|1|Axis Step
0071|SIEMENS SYNGO OBJECT GRAPHICS|51|SL|1|Axis Step Index
0071|SIEMENS SYNGO OBJECT GRAPHICS|52|CS|1|Axis Text Format
0071|SIEMENS SYNGO OBJECT GRAPHICS|53|CS|1|Axis Show Center Text Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|54|CS|1|Axis Show Tick Text Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|55|DS|3|Bitmap X Orientation
0071|SIEMENS SYNGO OBJECT GRAPHICS|56|DS|3|Bitmap Y Orientation
0071|SIEMENS SYNGO OBJECT GRAPHICS|57|OB|1|Graphic Blob
0071|SIEMENS SYNGO OBJECT GRAPHICS|58|CS|1|Graphic Interpolation
0071|SIEMENS SYNGO OBJECT GRAPHICS|59|DS|1|Graphic Angle
0071|SIEMENS SYNGO OBJECT GRAPHICS|60|DS|1|Graphic Size
0071|SIEMENS SYNGO OBJECT GRAPHICS|61|CS|1|Cut Line Side
0071|SIEMENS SYNGO OBJECT GRAPHICS|62|DS|1|Graphic Tip Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|63|DS|1|Cut Line Arrow Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|64|DS|1|Line Gap Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|65|DS|1|Graphic Circle Radius
0071|SIEMENS SYNGO OBJECT GRAPHICS|66|DS|1|Line Distance Move
0071|SIEMENS SYNGO OBJECT GRAPHICS|67|DS|1|Line Marker Length
0071|SIEMENS SYNGO OBJECT GRAPHICS|68|DS|3|Graphic Center
0071|SIEMENS SYNGO OBJECT GRAPHICS|69|DS|3|Range Center Area Top Left
0071|SIEMENS SYNGO OBJECT GRAPHICS|70|DS|3|Range Center Area Bottom Right
0071|SIEMENS SYNGO OBJECT GRAPHICS|71|DS|1|Range Tilt
0071|SIEMENS SYNGO OBJECT GRAPHICS|72|DS|1|Range Minimum Tilt
0071|SIEMENS SYNGO OBJECT GRAPHICS|73|DS|1|Range Maximum Tilt
0071|SIEMENS SYNGO OBJECT GRAPHICS|74|DS|1|Graphic Width
0071|SIEMENS SYNGO OBJECT GRAPHICS|75|DS|1|Range Minimum Width
0071|SIEMENS SYNGO OBJECT GRAPHICS|76|DS|1|Range Maximum Width
0071|SIEMENS SYNGO OBJECT GRAPHICS|77|DS|1|Graphic Height
0071|SIEMENS SYNGO OBJECT GRAPHICS|78|DS|1|Range Feed
0071|SIEMENS SYNGO OBJECT GRAPHICS|79|CS|1|Range Direction
0071|SIEMENS SYNGO OBJECT GRAPHICS|80|CS|1|Range Show Scans
0071|SIEMENS SYNGO OBJECT GRAPHICS|81|DS|1|Range Minimum Scan Distance
0071|SIEMENS SYNGO OBJECT GRAPHICS|82|CS|1|Range Orthogonal Height
0071|SIEMENS SYNGO OBJECT GRAPHICS|83|DS|3|Graphic Position
0071|SIEMENS SYNGO OBJECT GRAPHICS|84|CS|1|Graphic Closed Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|85|SL|1|Range Line Tip Mode
0071|SIEMENS SYNGO OBJECT GRAPHICS|86|SL|1|Graphic List Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|87|CS|1|Axis Flip Text Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|88|CS|1|Curve Diagram Type
0071|SIEMENS SYNGO OBJECT GRAPHICS|89|DS|1|Graphic Start Angle
0071|SIEMENS SYNGO OBJECT GRAPHICS|90|DS|1|Graphic End Angle
0071|SIEMENS SYNGO OBJECT GRAPHICS|91|IS|1|Live Wire Smoothness
0071|SIEMENS SYNGO OBJECT GRAPHICS|92|CS|1|Live Wire Spline Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|93|CS|1|Ellipse Circle Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|94|CS|1|Graphic Square Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|95|DS|1|Curve Section Start Index
0071|SIEMENS SYNGO OBJECT GRAPHICS|96|DS|1|Curve Section End Index
0071|SIEMENS SYNGO OBJECT GRAPHICS|97|DS|1|Marker Alpha
0071|SIEMENS SYNGO OBJECT GRAPHICS|98|IS|1|Table Row Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|99|IS|1|Table Column Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|9a|DS|1|Table Row Height
0071|SIEMENS SYNGO OBJECT GRAPHICS|9b|DS|1|Table Column Width
0071|SIEMENS SYNGO OBJECT GRAPHICS|9c|IS|1|Rectangle Selection Segment Offset
0071|SIEMENS SYNGO OBJECT GRAPHICS|9d|CS|1|Graphic Text
0071|SIEMENS SYNGO OBJECT GRAPHICS|a0|SL|1|Axis Tick Spacing Coordinate System
0071|SIEMENS SYNGO OBJECT GRAPHICS|a1|CS|1|Axis Diagram Grid Type
0071|SIEMENS SYNGO OBJECT GRAPHICS|a2|SL|1|Polar Plot Circle Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|a3|SL|1|Polar Plot Lines-per-Circle
0071|SIEMENS SYNGO OBJECT GRAPHICS|a4|SL|1|Polar Plot Compartment Count
0071|SIEMENS SYNGO OBJECT GRAPHICS|a5|SL|1|Polar Plot Radius Weight
0071|SIEMENS SYNGO OBJECT GRAPHICS|a6|DS|1|Circle Segment Outer Radius
0071|SIEMENS SYNGO OBJECT GRAPHICS|a7|CS|1|Circle Segment Clockwise Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|a8|CS|1|Axis Diagram Auto Resize Flag
0071|SIEMENS SYNGO OBJECT GRAPHICS|a9|DS|1|Axis Diagram Step Start
0071|SIEMENS SYNGO OBJECT GRAPHICS|b0|CS|1|Group Root
0071|SIEMENS SYNGO OBJECT GRAPHICS|b1|ST|1|Group Name
0071|SIEMENS SYNGO OBJECT GRAPHICS|b2|SQ|1|Graphic Annotation Sequence
0071|SIEMENS SYNGO OBJECT GRAPHICS|b3|SL|1|Text Minimum Height
0071|SIEMENS SYNGO OBJECT GRAPHICS|b4|DS|1|Text Font Scaling Factor
0071|SIEMENS SYNGO OBJECT GRAPHICS|b5|SL|2|Text Maximum Extensions
0071|SIEMENS SYNGO OBJECT GRAPHICS|b6|CS|1|Text Segment Size
0071|SIEMENS SYNGO OBJECT GRAPHICS|b7|SL|1|Graphic Object Reference Label
0073|SIEMENS SYNGO LAYOUT PROTOCOL|02|US|1|Hanging Protocol Excellence Rank
0073|SIEMENS SYNGO LAYOUT PROTOCOL|04|CS|1|Template Data Role ID
0073|SIEMENS SYNGO LAYOUT PROTOCOL|06|CS|1|Data Sharing Flag
0073|SIEMENS SYNGO LAYOUT PROTOCOL|08|SQ|1|Bagging Operations Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|10|LO|1|Synchronization Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|12|LO|1|Custom Filter Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|14|LO|1|Custom Sorter Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|16|CS|1|Reference Template Data Role ID
0073|SIEMENS SYNGO LAYOUT PROTOCOL|18|CS|1|Model Template Data Role ID
0073|SIEMENS SYNGO LAYOUT PROTOCOL|20|DT|1-n|Selector DT Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|22|DA|1-n|Selector DA Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|24|TM|1-n|Selector TM Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|26|UI|1-n|Selector UI Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|28|CS|1|Referenced Template Data Role
0073|SIEMENS SYNGO LAYOUT PROTOCOL|30|SQ|1|Custom Property Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|32|CS|1|Custom Property Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|34|LO|1|Custom Property Name
0073|SIEMENS SYNGO LAYOUT PROTOCOL|36|LO|1|Custom Property Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|38|SQ|1|Layout Property Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|40|SQ|1|Synchronization Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|42|CS|1|Presentation Creator Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|44|CS|1|Cine Navigation Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|48|LO|1|Semantic Naming Strategy
0073|SIEMENS SYNGO LAYOUT PROTOCOL|50|LO|1|Parameter String
0073|SIEMENS SYNGO LAYOUT PROTOCOL|52|CS|1|Sorting Order
0073|SIEMENS SYNGO LAYOUT PROTOCOL|54|CS|1|syngo Template Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|56|CS|1|Sorter Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|58|SH|1|Data Display Protocol Version
0073|SIEMENS SYNGO LAYOUT PROTOCOL|5a|CS|1|Timepoint Value
0073|SIEMENS SYNGO LAYOUT PROTOCOL|5b|CS|1|Sharing Group Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|5c|CS|1|Template Selector Operator
0073|SIEMENS SYNGO LAYOUT PROTOCOL|5d|CS|1|Sharing Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|60|SQ|1|Viewport Definitions Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|62|CS|1|Protocol Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|64|SQ|1|Template Selector Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|66|CS|1|Default Template
0073|SIEMENS SYNGO LAYOUT PROTOCOL|68|CS|1|Is Preferred
0073|SIEMENS SYNGO LAYOUT PROTOCOL|6a|SQ|1|Timepoint Initial Value Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|6c|CS|1|Timepoint Variable
0073|SIEMENS SYNGO LAYOUT PROTOCOL|70|SH|1|Display Protocol Name
0073|SIEMENS SYNGO LAYOUT PROTOCOL|72|LO|1|Display Protocol Description
0073|SIEMENS SYNGO LAYOUT PROTOCOL|74|CS|1|Display Protocol Level
0073|SIEMENS SYNGO LAYOUT PROTOCOL|76|LO|1|Display Protocol Creator
0073|SIEMENS SYNGO LAYOUT PROTOCOL|78|DT|1|Display Protocol Creation Datetime
0073|SIEMENS SYNGO LAYOUT PROTOCOL|7a|UI|1|Referenced Data Protocol
0073|SIEMENS SYNGO LAYOUT PROTOCOL|7c|US|1|Display Protocol Excellence Rank
0073|SIEMENS SYNGO LAYOUT PROTOCOL|7e|SQ|1|Layout Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|80|US|1|Layout Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|82|LO|1|Layout Description
0073|SIEMENS SYNGO LAYOUT PROTOCOL|84|SQ|1|Segment Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|86|US|1|Segment Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|88|LO|1|Segment Description
0073|SIEMENS SYNGO LAYOUT PROTOCOL|8a|CS|1|Segment Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|8c|US|1|Tile Horizontal Dimension
0073|SIEMENS SYNGO LAYOUT PROTOCOL|8e|US|1|Tile Vertical Dimension
0073|SIEMENS SYNGO LAYOUT PROTOCOL|90|CS|1|Fill Order
0073|SIEMENS SYNGO LAYOUT PROTOCOL|92|CS|1|Segment Small Scroll Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|94|US|1|Segment Small Scroll Amount
0073|SIEMENS SYNGO LAYOUT PROTOCOL|96|CS|1|Segment Large Scroll Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|98|US|1|Segment Large Scroll Amount
0073|SIEMENS SYNGO LAYOUT PROTOCOL|9a|US|1|Segment Overlap Priority
0073|SIEMENS SYNGO LAYOUT PROTOCOL|9c|SQ|1|Data Role View Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|9e|US|1|Data Role View Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|a2|US|1|Referenced Data Role
0073|SIEMENS SYNGO LAYOUT PROTOCOL|a4|CS|1|Sharing Enabled
0073|SIEMENS SYNGO LAYOUT PROTOCOL|a8|US|2-n|Referenced Data Role Views
0073|SIEMENS SYNGO LAYOUT PROTOCOL|b0|SH|1|Data Protocol Name
0073|SIEMENS SYNGO LAYOUT PROTOCOL|b2|LO|1|Data Protocol Description
0073|SIEMENS SYNGO LAYOUT PROTOCOL|b4|CS|1|Data Protocol Level
0073|SIEMENS SYNGO LAYOUT PROTOCOL|b6|LO|1|Data Protocol Creator
0073|SIEMENS SYNGO LAYOUT PROTOCOL|b8|DT|1|Data Protocol Creation Datetime
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ba|US|1|Data Protocol Excellence Rank
0073|SIEMENS SYNGO LAYOUT PROTOCOL|bc|SQ|1|Data Protocol Definition Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|be|SQ|1|Data Role Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|c0|US|1|Data Role Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|c2|SH|1|Data Role Name
0073|SIEMENS SYNGO LAYOUT PROTOCOL|c6|SQ|1|Selector Operations Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|c8|CS|1|Selector Usage Flag
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ca|CS|1|Select by Attribute Presence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|cc|CS|1|Select by Category
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ce|CS|1|Select by Operator
0073|SIEMENS SYNGO LAYOUT PROTOCOL|d0|LO|1|Custom Selector Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|d2|CS|1|Selector Operator
0073|SIEMENS SYNGO LAYOUT PROTOCOL|d4|CS|1|Reformatting Required
0073|SIEMENS SYNGO LAYOUT PROTOCOL|d6|SQ|1|Registration Data Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|d8|US|1|Reference Data Role Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|da|SQ|1|Model Data Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|dc|US|1|Model Data Role Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|de|SQ|1|Fusion Display Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|e0|FD|1|Transparency
0073|SIEMENS SYNGO LAYOUT PROTOCOL|e2|CS|1|Time Point
0073|SIEMENS SYNGO LAYOUT PROTOCOL|e4|LO|1|First Time Point Token
0073|SIEMENS SYNGO LAYOUT PROTOCOL|e6|LO|1|Last Time Point Token
0073|SIEMENS SYNGO LAYOUT PROTOCOL|e8|LO|1|Intermediate Time Point Token
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ea|SQ|1|Data Processor Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ec|LO|1|Data Processor Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ee|SQ|1|Template Data Role Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|f0|SQ|1|View Sequence
0073|SIEMENS SYNGO LAYOUT PROTOCOL|f4|LO|1|View Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|f6|LO|1|Custom Bagging Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|f8|US|1|Referenced Display Segment Number
0073|SIEMENS SYNGO LAYOUT PROTOCOL|fa|LO|1|Data Role Type
0073|SIEMENS SYNGO LAYOUT PROTOCOL|46|CS|1|Internal Flag
0073|SIEMENS SYNGO LAYOUT PROTOCOL|fc|CS|1|Unassigned Flag
0073|SIEMENS SYNGO LAYOUT PROTOCOL|fe|CS|1|Initial Display Scroll Position
0073|SIEMENS SYNGO LAYOUT PROTOCOL|ff|LO|1|VRT Preset
0091|SIENET|20|PN|1|RIS Patient Name
0093|SIENET|02|LO|1|Unknown
0095|SIENET|0c|SL|1|Unknown
0095|SIENET|20|PN|1|RIS Patient Name
0097|SIENET|03|SL|1|Unknown
0097|SIENET|05|LO|1|Unknown
0099|SIENET|05|SL|1|Unknown
00a5|SIENET|05|LO|1|Unknown
7fe3|SIEMENS MED NM|16|OW|1|Unknown
7fe3|SIEMENS MED NM|1b|OW|1|Unknown
7fe3|SIEMENS MED NM|1c|OW|1|Unknown
7fe3|SIEMENS MED NM|1e|OW|1|Unknown
7fe3|SIEMENS MED NM|26|OW|1|Unknown
7fe3|SIEMENS MED NM|27|OW|1|Unknown
7fe3|SIEMENS MED NM|28|OW|1|Unknown
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|10|LO|1|Evidence Document Template Name
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|11|DS|1|Evidence Document Template Version
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|20|OB|1|Clinical Finding Data
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|21|OB|1|Metadata
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|30|DS|1|Implementation Version
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|40|OB|1|Predecessor
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|50|LO|1|Logical ID
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|60|OB|1|Application Data
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|70|LO|1|Owner Clinical Task Name
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|71|LO|1|Owner Task Name
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|72|OB|1|Owner Supported Templates
0077|SIEMENS SYNGO EVIDENCE DOCUMENT DATA|80|OB|1|Volume Catalog
0021|syngoDynamics_Reporting|ad|OB|1|Data
0021|SIEMENS MR N3D|4a|SQ|1|Ortho MPR ColorLUT DR Sequence
0087|SIEMENS SYNGO ENCAPSULATED DOCUMENT DATA|20|OB|1|Study Model
0087|SIEMENS SYNGO ENCAPSULATED DOCUMENT DATA|30|OB|1|Report XML Schema
0087|SIEMENS SYNGO ENCAPSULATED DOCUMENT DATA|40|OB|1|Report Identifier
0029|SIEMENS SYNGO 3D FUSION MATRIX|08|UI|1|Object Series Instance UID
0029|SIEMENS SYNGO 3D FUSION MATRIX|09|UI|1|Model Series Instance UID
0029|SIEMENS SYNGO 3D FUSION MATRIX|10|UI|1|Matrix Referenced Series Instance UID
0019|SIEMENS Ultrasound SC2000|2d|US|1|B-mode Tint Index
0019|SIEMENS Ultrasound SC2000|72|US|1|Doppler Tint Index
0019|SIEMENS Ultrasound SC2000|88|US|1|M-mode Tint Index
0019|SIEMENS Ultrasound SC2000|89|LO|1|Unknown
0119|SIEMENS Ultrasound SC2000|00|LO|1|Acoustic Meta Information Version
0119|SIEMENS Ultrasound SC2000|01|UN|1|Common Acoustic Meta Information
0119|SIEMENS Ultrasound SC2000|02|SQ|1|Multi Stream Sequence
0119|SIEMENS Ultrasound SC2000|03|SQ|1|Acoustic Data Sequence
0119|SIEMENS Ultrasound SC2000|04|UN|1|Per Transaction Acoustic Control Information
0119|SIEMENS Ultrasound SC2000|05|UN|1|Acoustic Data Offset
0119|SIEMENS Ultrasound SC2000|06|UN|1|Acoustic Data Length
0119|SIEMENS Ultrasound SC2000|07|UN|1|Footer Offset
0119|SIEMENS Ultrasound SC2000|08|UN|1|Footer Length
0119|SIEMENS Ultrasound SC2000|09|UN|1|Acoustic Stream Number
0119|SIEMENS Ultrasound SC2000|10|UN|1|Acoustic Stream Type
0119|SIEMENS Ultrasound SC2000|11|UN|1|Stage Timer Time
0119|SIEMENS Ultrasound SC2000|12|UN|1|Stop Watch Time
0119|SIEMENS Ultrasound SC2000|13|UN|1|Volume Rate
0129|SIEMENS Ultrasound SC2000|00|SQ|1|MPR View Sequence
0129|SIEMENS Ultrasound SC2000|02|UI|1|Bookmark UID
0129|SIEMENS Ultrasound SC2000|03|UN|1|Plane Origin Vector
0129|SIEMENS Ultrasound SC2000|04|UN|1|Row Vector
0129|SIEMENS Ultrasound SC2000|05|UN|1|Column Vector
0129|SIEMENS Ultrasound SC2000|06|SQ|1|Visualization Sequence
0129|SIEMENS Ultrasound SC2000|07|UI|1|Bookmark UID
0129|SIEMENS Ultrasound SC2000|08|UN|1|Visualization Information
0129|SIEMENS Ultrasound SC2000|09|SQ|1|Application State Sequence
0129|SIEMENS Ultrasound SC2000|10|OB|1|Application State Information
0129|SIEMENS Ultrasound SC2000|11|SQ|1|Referenced Bookmark Sequence
0129|SIEMENS Ultrasound SC2000|12|UI|1|Referenced Bookmark UID
0129|SIEMENS Ultrasound SC2000|20|SQ|1|Cine Parameters Sequence
0129|SIEMENS Ultrasound SC2000|21|UN|1|Cine Parameters Schema
0129|SIEMENS Ultrasound SC2000|22|UN|1|Values of Cine Parameters
0129|SIEMENS Ultrasound SC2000|30|CS|1|Raw Data Object Type
0139|SIEMENS Ultrasound SC2000|01|SL|1|Physio Capture ROI
0149|SIEMENS Ultrasound SC2000|01|FD|1-n|Vector of BROI Points
0149|SIEMENS Ultrasound SC2000|02|FD|1-n|Start/End Timestamps of Strip Stream
0149|SIEMENS Ultrasound SC2000|03|FD|1-n|Timestamps of Visible R-waves
7fd1|SIEMENS Ultrasound SC2000|01|UN|1|Acoustic Image and Footer Data
7fd1|SIEMENS Ultrasound SC2000|09|UN|1|Volume Version ID
7fd1|SIEMENS Ultrasound SC2000|10|UN|1|Volume Payload
7fd1|SIEMENS Ultrasound SC2000|11|UN|1|After Payload
7fdf|SIEMENS SYNGO DATA PADDING|fc|OB|1|Pixel Data Leading Padding
0019|SIEMENS MR HEADER|08|CS|1|Unknown
0019|SIEMENS MR HEADER|09|LO|1|Unknown
0019|SIEMENS MR HEADER|0a|US|1|Number of Images in Mosaic
0019|SIEMENS MR HEADER|0b|DS|1|Slice Measurement Duration
0019|SIEMENS MR HEADER|0c|IS|1|B Value
0019|SIEMENS MR HEADER|0d|CS|1|Diffusion Directionality
0019|SIEMENS MR HEADER|0e|FD|3|Diffusion Gradient Direction
0019|SIEMENS MR HEADER|0f|SH|1|Gradient Mode
0019|SIEMENS MR HEADER|11|SH|1|Flow Compensation
0019|SIEMENS MR HEADER|12|SL|3|Table Position Origin
0019|SIEMENS MR HEADER|13|SL|3|Ima Abs Table Position
0019|SIEMENS MR HEADER|14|IS|3|Ima Rel Table Position
0019|SIEMENS MR HEADER|15|FD|3|Slice Position PCS
0019|SIEMENS MR HEADER|16|DS|1|Time After Start
0019|SIEMENS MR HEADER|17|DS|1|Slice Resolution
0019|SIEMENS MR HEADER|18|IS|1|Real Dwell Time
0019|SIEMENS MR HEADER|23|IS|1|Unknown
0019|SIEMENS MR HEADER|25|FD|1-n|Unknown
0019|SIEMENS MR HEADER|26|FD|1-n|Unknown
0019|SIEMENS MR HEADER|27|FD|6|B Matrix
0019|SIEMENS MR HEADER|28|FD|1|Bandwidth per Pixel Phase Encode
0019|SIEMENS MR HEADER|29|FD|1-n|Mosaic Ref Acq Times
0021|SIEMENS SERIES SHADOW ATTRIBUTES|01|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|02|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|03|OB|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|04|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|05|IS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|06|LO|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|07|LO|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|08|SH|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|09|LO|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|0a|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|0c|SH|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|0d|US|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|0f|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|10|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|11|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|12|FD|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|13|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|14|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|16|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|17|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|18|SH|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|19|OB|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|1a|LO|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|1b|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|1c|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|1d|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|1f|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|22|SH|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|23|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|25|SL|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|26|IS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|27|US|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2a|IS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2b|ST|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2c|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2d|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2e|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|2f|DS|1-n|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|30|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|31|IS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|32|SS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|33|SH|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|34|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|35|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|36|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|38|DS|1|Unknown
0021|SIEMENS SERIES SHADOW ATTRIBUTES|3b|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|01|US|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|02|FD|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|03|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|04|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|05|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|06|LO|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|1a|SH|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|1c|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|1f|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|20|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|22|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|24|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|25|LT|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|26|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|27|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|2a|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|2b|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|2c|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|2d|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|2e|UL|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|33|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|34|FD|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|35|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|37|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|3a|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|3b|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|3c|FD|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|3d|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|3f|SH|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|40|DS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|41|SH|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|42|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|43|LT|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|44|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|45|SL|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|46|FD|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|47|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|48|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|49|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|4b|LT|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|4e|IS|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|4f|LO|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|51|UL|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|52|US|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|53|FD|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|54|US|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|56|LO|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|58|SH|1|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|59|IS|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|5a|FD|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|5b|FD|1-n|Unknown
0021|SIEMENS IMAGE SHADOW ATTRIBUTES|5e|IS|1|Unknown
0021|SIEMENS MR IMA|01|SQ|1|MR Image Sequence
0021|SIEMENS MR N3D|30|SQ|1|Background Color DR Sequence
0021|SIEMENS MR N3D|31|DS|3|Background Color
0021|SIEMENS MR N3D|36|SQ|1|Field Map DR Sequence
0021|SIEMENS MR N3D|37|CS|1|Visible
0021|SIEMENS MR N3D|38|DS|3|Tinting Color
0021|SIEMENS MR N3D|39|CS|1|Tinting Enabled
0021|SIEMENS MR N3D|3a|LO|1|Volume ID
0021|SIEMENS MR N3D|3b|LO|1|Volume ID As Bound
0021|SIEMENS MR N3D|41|SQ|1|Floating MPR Color LUT DR Sequence
0021|SIEMENS MR N3D|42|DS|1|RGBA LUT
0021|SIEMENS MR N3D|43|DS|1|Blend Factor
0021|SIEMENS MR N3D|44|SQ|1|RGBA LUT Data Sequence
0021|SIEMENS MR N3D|45|OB|1|Color LUT
0021|SIEMENS MR N3D|4b|SQ|1|VRT Color LUT DR Sequence
0021|SIEMENS MR N3D|4d|SQ|1|Pwl Transfer Function Data Sequence
0021|SIEMENS MR N3D|4c|SQ|1|Pwl Transfer Function Sequence
0021|SIEMENS MR N3D|4e|DS|1|Pwl Vertex Index
0021|SIEMENS MR N3D|50|SQ|1|Pwl Vertex Sequence
0021|SIEMENS MR N3D|51|SQ|1|Floating MPR Render DR Sequence
0021|SIEMENS MR N3D|52|CS|1|Primary Show Hide
0021|SIEMENS MR N3D|56|CS|1|Alpha Dependent Fieldmap
0021|SIEMENS MR N3D|57|LO|1|Volume Filter
0021|SIEMENS MR N3D|5a|SQ|1|Ortho MPR Render DR Sequence
0021|SIEMENS MR N3D|5b|SQ|1|VRT Render DR Sequence
0021|SIEMENS MR N3D|53|CS|1|Secondary Show Hide
0021|SIEMENS MR N3D|54|LO|1|Primary Shading Index
0021|SIEMENS MR N3D|55|LO|1|Secondary Shading Index
0021|SIEMENS MR N3D|58|DS|3|Bounding Box Color
0021|SIEMENS MR N3D|59|CS|1|Scene Interaction On
0021|SIEMENS MR N3D|60|SQ|6|Clip Plane DR Sequence
0021|SIEMENS MR N3D|61|DS|3|Plane Center
0021|SIEMENS MR N3D|62|DS|3|Plane Normal
0021|SIEMENS MR N3D|63|DS|2|Plane Scale
0021|SIEMENS MR N3D|64|CS|1|Plane Enable GL Clip
0021|SIEMENS MR N3D|65|DS|1|Plane Handle Ratio
0021|SIEMENS MR N3D|66|DS|24|Plane Bounding Points
0021|SIEMENS MR N3D|67|DS|16|Plane Motion Matrix
0021|SIEMENS MR N3D|68|DS|1|Plane Shift Velocity
0021|SIEMENS MR N3D|69|CS|1|Plane Enabled
0021|SIEMENS MR N3D|6a|DS|1|Plane Rotate Velocity
0021|SIEMENS MR N3D|6b|CS|1|Plane Show Graphics
0021|SIEMENS MR N3D|73|CS|1|Plane Single Selection Mode
0021|SIEMENS MR N3D|74|CS|1|Plane Alignment
0021|SIEMENS MR N3D|75|CS|1|Plane Selected
0021|SIEMENS MR N3D|70|SQ|1|Split Plane DR Sequence
0021|SIEMENS MR N3D|71|SQ|3|Floating MPR DR Sequence
0021|SIEMENS MR N3D|6e|CS|1|Plane MPR Locked
0021|SIEMENS MR N3D|6f|CS|1|Plane Scaling Disabled
0021|SIEMENS MR N3D|72|SQ|3|Ortho MPR DR Sequence
0021|SIEMENS MR N3D|6c|DS|1|Offset
0021|SIEMENS MR N3D|6d|CS|1|Ortho MPR At Bounding Box
0021|SIEMENS MR N3D|76|SQ|1|Clustering DR Sequence
0021|SIEMENS MR N3D|77|DS|1|Cluster Size
0021|SIEMENS MR N3D|78|CS|1|Clustering Enabled
0021|SIEMENS MR N3D|79|LO|1|Cluster Mask Vol ID
0021|SIEMENS MR N3D|80|SQ|1|Head Masking DR Sequence
0021|SIEMENS MR N3D|81|DS|2|Masking Range
0021|SIEMENS MR N3D|82|CS|1|Mask Enabled
0021|SIEMENS MR N3D|83|SQ|1|Brain Masking DR Sequence
0021|SIEMENS MR N3D|84|SQ|1|Masking Status DR Sequence
0021|SIEMENS MR N3D|85|SQ|1|VRT Masking DR Sequence
0021|SIEMENS MR N3D|86|SQ|1|Ortho MPR Masking DR Sequence
0021|SIEMENS MR N3D|87|SQ|1|Floating MPR Masking DR Sequence
0021|SIEMENS MR N3D|88|SQ|1|Align DR Sequence
0021|SIEMENS MR N3D|89|DS|16|Registration Matrix
0021|SIEMENS MR N3D|90|SQ|1|Functional Evaluation DR Sequence
0021|SIEMENS MR N3D|91|DS|1-n|Frame Acquition Numbers
0021|SIEMENS MR N3D|92|CS|1|Show Cursor
0021|SIEMENS MR N3D|93|DS|1|Current Frame
0021|SIEMENS MR N3D|94|DS|1-n|Plot Area
0021|SIEMENS MR N3D|95|DS|2|Plot Text Position
0021|SIEMENS MR N3D|96|DS|1-n|Base Line Points
0021|SIEMENS MR N3D|97|DS|1-n|Active Points
0021|SIEMENS MR N3D|98|CS|1|Show Label
0021|SIEMENS MR N3D|99|CS|1|Mean Plot
0021|SIEMENS MR N3D|9a|CS|1|Motion Plot
0021|SIEMENS MR N3D|9b|CS|1|Activate Normallized Curve
0021|SIEMENS MR N3D|9c|DS|1|Plot Size
0021|SIEMENS MR N3D|a0|SQ|4|PlotDR Sequence
0021|SIEMENS MR N3D|a1|LO|1|Title
0021|SIEMENS MR N3D|a2|CS|1|Auto Scale
0021|SIEMENS MR N3D|a3|DS|1|Fixed Scale
0021|SIEMENS MR N3D|a4|DS|3|Background Color
0021|SIEMENS MR N3D|a5|LO|1|Label X
0021|SIEMENS MR N3D|a6|LO|1|Label Y
0021|SIEMENS MR N3D|a7|CS|1|Legend
0021|SIEMENS MR N3D|a8|CS|1|Scroll Bar X
0021|SIEMENS MR N3D|a9|CS|1|Scroll Bar Y
0021|SIEMENS MR N3D|aa|LO|1|Connect Scroll X
0021|SIEMENS MR N3D|ab|LO|1|Plot ID
0021|SIEMENS MR N3D|ac|DS|1|Plot Position
0021|SIEMENS MR N3D|b0|SQ|1|Curve DR Sequence
0021|SIEMENS MR N3D|b1|LO|1|Curve ID
0021|SIEMENS MR N3D|b2|LO|1|Plot Type
0021|SIEMENS MR N3D|b3|DS|1-n|Curve Values
0021|SIEMENS MR N3D|b4|DS|3|Line Color
0021|SIEMENS MR N3D|b5|DS|3|Marker Color
0021|SIEMENS MR N3D|b6|CS|1|Line Filled
0021|SIEMENS MR N3D|b7|LO|1|Label
0021|SIEMENS MR N3D|b8|CS|1|Show Marker
0021|SIEMENS MR N3D|b9|LO|1|Marker Shape
0021|SIEMENS MR N3D|ba|LO|1|Smoothing Algo
0021|SIEMENS MR N3D|bb|DS|1|Marker Size
0021|SIEMENS MR N3D|bc|LO|1|Line Style
0021|SIEMENS MR N3D|bd|LO|1|Line Pattern
0021|SIEMENS MR N3D|be|DS|1|Line Width
0021|SIEMENS MR N3D|c0|SQ|1|VRT Filter DR Sequence
0021|SIEMENS MR N3D|c1|LO|1|Filter Type
0021|SIEMENS MR N3D|c2|CS|1|Current Active Plane
0021|SIEMENS MR PHOENIX ATTRIBUTES|01|UL|1|Mds Mode Mask
0021|SIEMENS MR PHOENIX ATTRIBUTES|02|US|1|Dixon
0021|SIEMENS MR PHOENIX ATTRIBUTES|03|LT|1|Sequence File Name
0021|SIEMENS MR PHOENIX ATTRIBUTES|f1|UL|1|Count of Pseudo Attributes
0021|SIEMENS MR SDS 01|fe|SQ|1|Siemens MR SDS Sequence
0021|SIEMENS MR SDS 01|01|IS|1|Used Patient Weight
0021|SIEMENS MR SDS 01|02|DS|3|SAR Whole Body
0021|SIEMENS MR SDS 01|03|OB|1|MR Protocol
0021|SIEMENS MR SDS 01|04|DS|1|Slice Array Concatenations
0021|SIEMENS MR SDS 01|05|IS|3|Rel Table Position
0021|SIEMENS MR SDS 01|06|LO|1|Coil For Gradient
0021|SIEMENS MR SDS 01|07|LO|1|Long Model Name
0021|SIEMENS MR SDS 01|08|SH|1|Gradient Mode
0021|SIEMENS MR SDS 01|09|LO|1|PAT Mode Text
0021|SIEMENS MR SDS 01|0a|DS|1|SW Correction Factor
0021|SIEMENS MR SDS 01|0b|DS|1|RF Power Error Indicator
0021|SIEMENS MR SDS 01|0c|SH|1|Positive PCS Directions
0021|SIEMENS MR SDS 01|0d|US|1|Protocol Change History
0021|SIEMENS MR SDS 01|0e|LO|1|Data File Name
0021|SIEMENS MR SDS 01|0f|DS|3|Stimlim
0021|SIEMENS MR SDS 01|10|IS|1|MR Protocol Version
0021|SIEMENS MR SDS 01|11|DS|1|Phase Gradient Amplitude
0021|SIEMENS MR SDS 01|12|FD|1|Readout OS
0021|SIEMENS MR SDS 01|13|DS|1|tpuls max
0021|SIEMENS MR SDS 01|14|IS|1|Number of Prescans
0021|SIEMENS MR SDS 01|15|FL|1|Measurement Index
0021|SIEMENS MR SDS 01|16|DS|1|dBdt Threshold
0021|SIEMENS MR SDS 01|17|DS|1|Selection Gradient Amplitude
0021|SIEMENS MR SDS 01|18|SH|1|RF SWD Most Critical Aspect
0021|SIEMENS MR SDS 01|19|OB|1|MR Phoenix Protocol
0021|SIEMENS MR SDS 01|1a|LO|1|Coil String
0021|SIEMENS MR SDS 01|1b|DS|1|Slice Resolution
0021|SIEMENS MR SDS 01|1c|DS|3|Stim max online
0021|SIEMENS MR SDS 01|1d|IS|1|Operation Mode Flag
0021|SIEMENS MR SDS 01|1e|FL|16|Auto Align Matrix
0021|SIEMENS MR SDS 01|1f|DS|2|Coil Tuning Reflection
0021|SIEMENS MR SDS 01|20|UI|1|Representative Image
0021|SIEMENS MR SDS 01|22|SH|1|Sequence File Owner
0021|SIEMENS MR SDS 01|23|IS|1|RF Watchdog Mask
0021|SIEMENS MR SDS 01|24|LO|1|Post Proc Protocol
0021|SIEMENS MR SDS 01|25|SL|3|Table Position Origin
0021|SIEMENS MR SDS 01|26|IS|32|Misc Sequence Param
0021|SIEMENS MR SDS 01|27|US|1|Isocentered
0021|SIEMENS MR SDS 01|2a|IS|1-n|Coil ID
0021|SIEMENS MR SDS 01|2b|ST|1|Pat Rein Pattern
0021|SIEMENS MR SDS 01|2c|DS|3|SED
0021|SIEMENS MR SDS 01|2d|DS|3|SAR Most Critical Aspect
0021|SIEMENS MR SDS 01|2e|IS|1|Stimm on mode
0021|SIEMENS MR SDS 01|2f|DS|3|Gradient Delay Time
0021|SIEMENS MR SDS 01|30|DS|1|Readout Gradient Amplitude
0021|SIEMENS MR SDS 01|31|IS|1|Abs Table Position
0021|SIEMENS MR SDS 01|32|SS|1|RF SWD Operation Mode
0021|SIEMENS MR SDS 01|33|SH|1|Coil for Gradient2
0021|SIEMENS MR SDS 01|34|DS|1|Stim Factor
0021|SIEMENS MR SDS 01|35|DS|1|Stim max ges norm online
0021|SIEMENS MR SDS 01|36|DS|1|dBdt max
0021|SIEMENS MR SDS 01|38|DS|1|Transmitter Calibration
0021|SIEMENS MR SDS 01|39|OB|1|MR EVA Protocol
0021|SIEMENS MR SDS 01|3b|DS|1|dBdt Limit
0021|SIEMENS MR SDS 01|3c|OB|1|VF Model Info
0021|SIEMENS MR SDS 01|3d|CS|1|Phase Slice Oversampling
0021|SIEMENS MR SDS 01|3e|OB|1|VF Settings
0021|SIEMENS MR SDS 01|3f|UT|1|Auto Align Data
0021|SIEMENS MR SDS 01|40|UT|1|FMRI Model Parameters
0021|SIEMENS MR SDS 01|41|UT|1|FMRI Model Info
0021|SIEMENS MR SDS 01|42|UT|1|FMRI External Parameters
0021|SIEMENS MR SDS 01|43|UT|1|FMRI External Info
0021|SIEMENS MR SDS 01|44|DS|2|B1 RMS
0021|SIEMENS MR SDS 01|45|CS|1|B1 RMS Supervision
0021|SIEMENS MR SDS 01|46|DS|1|Tales Reference Power
0021|SIEMENS MR SDS 01|47|CS|1|Safety Standard
0021|SIEMENS MR SDS 01|48|CS|1|DICOM Image Flavor
0021|SIEMENS MR SDS 01|49|CS|1|DICOM Acquisition Contrast
0021|SIEMENS MR SDS 01|50|US|1|RF Echo Train Length 4MF
0021|SIEMENS MR SDS 01|51|US|1|Gradient Echo Train Length 4MF
0021|SIEMENS MR SDS 01|52|LO|1|Version Info
0021|SIEMENS MR SDS 01|53|CS|1|Laterality 4MF
0021|SIEMENS MR MRS 05|01|FD|1|Transmitter Reference Amplitude
0021|SIEMENS MR MRS 05|02|US|1|Hamming Filter Width
0021|SIEMENS MR MRS 05|03|FD|3|CSI Gridshift Vector
0021|SIEMENS MR MRS 05|04|FD|1|Mixing Time
0021|SIEMENS MR MRS 05|40|CS|1|Series Protocol Instance
0021|SIEMENS MR MRS 05|41|CS|1|Spectro Result Type
0021|SIEMENS MR MRS 05|42|CS|1|Spectro Result Extend Type
0021|SIEMENS MR MRS 05|43|CS|1|Post Proc Protocol
0021|SIEMENS MR MRS 05|44|CS|1|Rescan Level
0021|SIEMENS MR MRS 05|45|OF|1|Spectro Algo Result
0021|SIEMENS MR MRS 05|46|OF|1|Spectro Display Params
0021|SIEMENS MR MRS 05|47|IS|1|Voxel Number
0021|SIEMENS MR MRS 05|48|SQ|1|APR Sequence
0021|SIEMENS MR MRS 05|49|CS|1|Sync Data
0021|SIEMENS MR MRS 05|4a|CS|1|Post Proc Detailed Protocol
0021|SIEMENS MR MRS 05|4b|CS|1|Spectro Result Extend Type Detailed
0025|SIEMENS MR EXTRACTED CSA HEADER|01|SQ|1|Extracted MR Header Information Sequence
0025|SIEMENS MR EXTRACTED CSA HEADER|02|LO|1|Extracted MR Header Creator Identification Code
0025|SIEMENS MR EXTRACTED CSA HEADER|03|AT|1|Extracted MR Header Tag
0051|SIEMENS MR HEADER|08|CS|1|CSA Image Header Type
0051|SIEMENS MR HEADER|09|LO|1|CSA Image Header Version
0051|SIEMENS MR HEADER|0a|LO|1|Unknown
0051|SIEMENS MR HEADER|0b|SH|1|Acquisition Matrix Text
0051|SIEMENS MR HEADER|0c|LO|1|Unknown
0051|SIEMENS MR HEADER|0d|SH|1|Unknown
0051|SIEMENS MR HEADER|0e|LO|1|Unknown
0051|SIEMENS MR HEADER|0f|LO|1|Coil String
0051|SIEMENS MR HEADER|11|LO|1|Unknown
0051|SIEMENS MR HEADER|12|SH|1|Unknown
0051|SIEMENS MR HEADER|13|SH|1|Positive PCS Directions
0051|SIEMENS MR HEADER|15|SH|1|Unknown
0051|SIEMENS MR HEADER|16|LO|1|Unknown
0051|SIEMENS MR HEADER|17|SH|1|Unknown
0051|SIEMENS MR HEADER|18|SH|1|Unknown
0051|SIEMENS MR HEADER|19|LO|1|Unknown
0021|SIEMENS MR SDI 02|01|US|1|Number of Images in Mosaic
0021|SIEMENS MR SDI 02|02|FD|3|Slice Normal Vector
0021|SIEMENS MR SDI 02|03|DS|1|Slice Measurement Duration
0021|SIEMENS MR SDI 02|04|DS|1|Time After Start
0021|SIEMENS MR SDI 02|05|IS|1|B Value
0021|SIEMENS MR SDI 02|06|LO|1|ICE Dims
0021|SIEMENS MR SDI 02|1a|SH|1|RF SWD Data Type
0021|SIEMENS MR SDI 02|1b|US|1|MoCoQ Measure
0021|SIEMENS MR SDI 02|1c|IS|1|Phase Encoding Direction Positive
0021|SIEMENS MR SDI 02|1d|OB|1|Pixel File
0021|SIEMENS MR SDI 02|1f|IS|1|FMRI Stimul Info
0021|SIEMENS MR SDI 02|20|DS|1|Voxel in Plane Rot
0021|SIEMENS MR SDI 02|21|CS|1|Diffusion Directionality 4MF
0021|SIEMENS MR SDI 02|22|DS|1|Voxel Thickness
0021|SIEMENS MR SDI 02|23|FD|6|B Matrix
0021|SIEMENS MR SDI 02|24|IS|1|Multistep Index
0021|SIEMENS MR SDI 02|25|LT|1|Comp Adjusted Param
0021|SIEMENS MR SDI 02|26|IS|1|Comp Algorithm
0021|SIEMENS MR SDI 02|27|DS|1|Voxel NormalC or
0021|SIEMENS MR SDI 02|29|SH|1|Flow Encoding Direction String
0021|SIEMENS MR SDI 02|2a|DS|1|Voxel Normal Sag
0021|SIEMENS MR SDI 02|2b|DS|1|Voxel Position Sag
0021|SIEMENS MR SDI 02|2c|DS|1|Voxel Normal Tra
0021|SIEMENS MR SDI 02|2d|DS|1|Voxel Position Tra
0021|SIEMENS MR SDI 02|2e|UL|1|Used Channel Mask
0021|SIEMENS MR SDI 02|2f|DS|1|Repetition Time Effective
0021|SIEMENS MR SDI 02|30|DS|6|CSI Image Orientation Patient
0021|SIEMENS MR SDI 02|32|DS|1|CSI Slice Location
0021|SIEMENS MR SDI 02|33|IS|1|Echo Column Position
0021|SIEMENS MR SDI 02|34|FD|1|Flow VENC
0021|SIEMENS MR SDI 02|35|IS|1|Measured Fourier Lines
0021|SIEMENS MR SDI 02|36|SH|1|LQ Algorithm
0021|SIEMENS MR SDI 02|37|DS|1|Voxel Position Cor
0021|SIEMENS MR SDI 02|38|IS|1|Filter2
0021|SIEMENS MR SDI 02|39|FD|1|FMRI Stimul Level
0021|SIEMENS MR SDI 02|3a|DS|1|Voxel Readout FOV
0021|SIEMENS MR SDI 02|3b|IS|1|Normalize Manipulated
0021|SIEMENS MR SDI 02|3c|FD|3|RBMoCoRot
0021|SIEMENS MR SDI 02|3d|IS|1|Comp Manual Adjusted
0021|SIEMENS MR SDI 02|3f|SH|1|Spectrum Text Region Label
0021|SIEMENS MR SDI 02|40|DS|1|Voxel Phase FOV
0021|SIEMENS MR SDI 02|41|SH|1|GSWD Data Type
0021|SIEMENS MR SDI 02|42|IS|1|Real Dwell Time
0021|SIEMENS MR SDI 02|43|LT|1|Comp Job ID
0021|SIEMENS MR SDI 02|44|IS|1|Comp Blended
0021|SIEMENS MR SDI 02|45|SL|3|Ima Abs Table Position
0021|SIEMENS MR SDI 02|46|FD|3|Diffusion Gradient Direction
0021|SIEMENS MR SDI 02|47|IS|1|Flow Encoding Direction
0021|SIEMENS MR SDI 02|48|IS|1|Echo Partition Position
0021|SIEMENS MR SDI 02|49|IS|1|Echo Line Position
0021|SIEMENS MR SDI 02|4b|LT|1|Comp Auto Param
0021|SIEMENS MR SDI 02|4c|IS|1|Original Image Number
0021|SIEMENS MR SDI 02|4d|IS|1|Original Series Number
0021|SIEMENS MR SDI 02|4e|IS|1|Actual 3D Ima Part Number
0021|SIEMENS MR SDI 02|4f|LO|1|Ima Coil String
0021|SIEMENS MR SDI 02|50|DS|2|CSI Pixel Spacing
0021|SIEMENS MR SDI 02|51|UL|1|Sequence Mask
0021|SIEMENS MR SDI 02|52|US|1|Image Group
0021|SIEMENS MR SDI 02|53|FD|1|Bandwidth Per Pixel Phase Encode
0021|SIEMENS MR SDI 02|54|US|1|Non Planar Image
0021|SIEMENS MR SDI 02|55|OB|1|Pixel File Name
0021|SIEMENS MR SDI 02|56|LO|1|Ima PAT Mode Text
0021|SIEMENS MR SDI 02|57|DS|3|CSI Image Position Patient
0021|SIEMENS MR SDI 02|58|SH|1|Acquisition Matrix Text
0021|SIEMENS MR SDI 02|59|IS|3|Ima Rel Table Position
0021|SIEMENS MR SDI 02|5a|FD|3|RBMoCoTrans
0021|SIEMENS MR SDI 02|5b|FD|3|Slice Position PCS
0021|SIEMENS MR SDI 02|5c|DS|1|CSI Slice Thickness
0021|SIEMENS MR SDI 02|5e|IS|1|Protocol Slice Number
0021|SIEMENS MR SDI 02|5f|IS|1|Filter1
0021|SIEMENS MR SDI 02|60|SH|1|Transmitting Coil
0021|SIEMENS MR SDI 02|61|DS|1|Number of Averages N4
0021|SIEMENS MR SDI 02|62|FD|1-n|Mosaic Ref Acq Times
0021|SIEMENS MR SDI 02|63|IS|1|Auto Inline Image Filter Enabled
0021|SIEMENS MR SDI 02|65|FD|1-n|QC Data
0021|SIEMENS MR SDI 02|66|LT|1|Exam Landmarks
0021|SIEMENS MR SDI 02|67|ST|1|Exam Data Role
0021|SIEMENS MR SDI 02|68|OB|1|MR Diffusion
0021|SIEMENS MR SDI 02|69|OB|1|Real World Value Mapping
0021|SIEMENS MR SDI 02|70|OB|1|Data Set Info
0021|SIEMENS MR SDI 02|71|UT|1|Used Channel String
0021|SIEMENS MR SDI 02|72|CS|1|Phase ContrastN4
0021|SIEMENS MR SDI 02|73|UT|1|MR Velocity Encoding
0021|SIEMENS MR SDI 02|74|FD|3|Velocity Encoding Direction N4
0021|SIEMENS MR SDI 02|75|CS|1-n|Image Type 4MF
0021|SIEMENS MR SDI 02|76|LO|1-n|Image History
0021|SIEMENS MR SDI 02|77|LO|1|SequenceI nfo
0021|SIEMENS MR SDI 02|78|CS|1-n|Image Type Visible
0021|SIEMENS MR SDI 02|79|CS|1|Distortion Correction Type
0021|SIEMENS MR SDI 02|80|CS|1|Image Filter Type
0021|SIEMENS MR SDI 02|fe|SQ|1|Siemens MR SDI Sequence
0021|SIEMENS MR CM 03|01|IS|1|Unknown
0021|SIEMENS MR CM 03|02|CS|1|Unknown
0021|SIEMENS MR PS 04|01|FD|1-n|Unknown
0021|SIEMENS MR FOR 06|01|LO|1|Unknown
0029|SIEMENS CT APPL DATASET|00|LT|1|Dual Energy Algorithm Parameters
0029|SIEMENS CT APPL DATASET|01|US|1|Valid CT Volume MBox Tasks
0029|SIEMENS CT APPL DATASET|02|LT|1|Scan Options
0029|SIEMENS CT APPL DATASET|03|ST|1|Acquisition Date and Time
0029|SIEMENS CT APPL DATASET|04|ST|1|Acquisition Number
0029|SIEMENS CT APPL DATASET|05|ST|1|Dynamic Data
0029|SIEMENS CT APPL DATASET|06|DS|6|Image Orientation Patient
0029|SIEMENS CT APPL DATASET|07|LT|1|Frame Of Reference Uid
0029|SIEMENS CT APPL DATASET|08|LT|1|Patient Position
0029|SIEMENS CT APPL DATASET|09|LT|1|Convolution Kernel
0029|SIEMENS CT APPL DATASET|10|LT|1|Kvp
0029|SIEMENS CT APPL DATASET|11|LT|1|Reconstruction Diameter
0029|SIEMENS CT APPL DATASET|12|LT|1|Rescale Intercept
0029|SIEMENS CT APPL DATASET|13|LT|1|Rescale Slope
0029|SIEMENS CT APPL DATASET|14|LT|1|Slice Thickness
0029|SIEMENS CT APPL DATASET|15|LT|1|Table Height
0029|SIEMENS CT APPL DATASET|16|LT|1|Gantry Detector Tilt
0029|SIEMENS CT APPL DATASET|17|LT|1|Pixel Spacing
0029|SIEMENS CT APPL DATASET|18|ST|1|Volume PatientPosition Not Equal
0029|SIEMENS CT APPL DATASET|19|ST|1|Volume LossyImageCompression Not Equal
0029|SIEMENS CT APPL DATASET|20|ST|1|Volume ConvolutionKernel Not Equal
0029|SIEMENS CT APPL DATASET|21|ST|1|Volume PixelSpacing Not Equal
0029|SIEMENS CT APPL DATASET|22|ST|1|Volume Kvp Not Equal
0029|SIEMENS CT APPL DATASET|23|ST|1|Volume ReconstructionDiameter Not Equal
0029|SIEMENS CT APPL DATASET|24|ST|1|Volume TableHeight Not Equal
0029|SIEMENS CT APPL DATASET|25|ST|1|Volume Has Gaps
0029|SIEMENS CT APPL DATASET|26|ST|1|Volume Number Of Missing Images
0029|SIEMENS CT APPL DATASET|27|ST|1|Volume Max Gap
0029|SIEMENS CT APPL DATASET|28|LT|1|Volume Position Of Gaps
0029|SIEMENS CT APPL DATASET|29|FD|1|Calibration Factor
0029|SIEMENS CT APPL DATASET|2a|CS|1|Flash Mode
0029|SIEMENS CT APPL DATASET|2b|LT|1|Warnings
0029|SIEMENS CT APPL DATASET|2c|ST|1|Volume HighBit Not Equal
0029|SIEMENS CT APPL DATASET|2d|ST|1|Volume ImageType Not Equal
0029|SIEMENS CT APPL DATASET|2e|ST|1|ImageType 0
0029|SIEMENS CT APPL DATASET|2f|ST|1|ImageType 1
0029|SIEMENS CT APPL DATASET|30|ST|1|ImageType 2
0029|SIEMENS CT APPL DATASET|31|ST|1|ImageType 3
0029|SIEMENS CT APPL DATASET|32|ST|1|PhotometricInterpretation not MONOCHROME2
0029|SIEMENS CT APPL DATASET|33|DA|1|First Acquisition Date
0029|SIEMENS CT APPL DATASET|34|DA|1|Last Acquisition Date
0029|SIEMENS CT APPL DATASET|35|TM|1|First Acquisition Time
0029|SIEMENS CT APPL DATASET|36|TM|1|Last Acquisition Time
0029|SIEMENS CT APPL DATASET|37|ST|1|Internal Data
0029|SIEMENS CT APPL DATASET|38|ST|1|Ranges SOM7
0029|SIEMENS CT APPL DATASET|39|LT|1|Calculated Gantry Detector Tilt
0029|SIEMENS CT APPL DATASET|40|ST|1|Volume Slice Distance
0029|SIEMENS CT APPL DATASET|41|DS|1|First Slice Z Coordinate 
0029|SIEMENS CT APPL DATASET|42|DS|1|Last Slice Z Coordinate 
0029|SIEMENS CT APPL DATASET|43|DS|1|Content DateTime
0029|SIEMENS CT APPL DATASET|44|DS|1|Delta Time
0029|SIEMENS CT APPL DATASET|45|DS|1|Frame Count
0029|SIEMENS CT APPL EVIDENCEDOCUMENT|00|UT|1|Private Task Datamodel
0029|SIEMENS CT APPL MEASUREMENT|00|UT|1|Oncology Segmentation Measurement Values
0029|SIEMENS CT APPL MEASUREMENT|01|ST|1|Oncology Measurement Recist Standard
0029|SIEMENS CT APPL MEASUREMENT|10|CS|1|DualEnergy ROI Annotation Mode
0029|SIEMENS CT APPL PRESENTATION|00|US|1|Translucent Mode
0029|SIEMENS CT APPL PRESENTATION|01|FD|1|Translucent Window Size
0029|SIEMENS CT APPL PRESENTATION|02|US|1|Panoramic Mode
0029|SIEMENS CT APPL PRESENTATION|03|FD|1|Panoramic Inner Width
0029|SIEMENS CT APPL PRESENTATION|04|US|1|Display Unseen Areas
0029|SIEMENS CT APPL PRESENTATION|05|US|4|Unseen Areas Color
0029|SIEMENS CT APPL PRESENTATION|06|US|1|Display Tagged Data
0029|SIEMENS CT APPL PRESENTATION|07|US|4|Tagged Color
0029|SIEMENS CT APPL PRESENTATION|08|UL|1|Tagged Sample Thickness
0029|SIEMENS CT APPL PRESENTATION|09|SL|1|Tagged Threshold
0029|SIEMENS CT APPL PRESENTATION|10|US|1|Kernel Filter
0029|SIEMENS CT APPL TMP DATAMODEL|00|OB|1|CT Task Common DataModel
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|00|UN|1|Release Version
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|03|UN|1|Volume Acquisition Duration
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|04|UN|1|Volume Raw Data Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|05|UN|1|Scan Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|06|UN|1|Z Lateral Min
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|07|UN|1|Z Lateral Span
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|08|UN|1|Z Radius of Curvature
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|09|UN|1|Wobble Correction
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|10|UN|1|Scale Along Width
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|11|UN|1|Scale Along Height
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|12|UN|1|Scale Along Depth
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|13|UN|1|Buffer Size
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|14|UN|1|Acquisition Rate
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|15|UN|1|Depth Min cm
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|16|UN|1|Is Left Right Flipped Enabled
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|17|UN|1|Is Up Down Flipped Enabled
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|18|UN|1|Is Volume Geom Accurate
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|19|UN|1|BByte Mask Offset
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|20|UN|1|BByte Mask Size
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|22|UN|1|Acq Plane Rotation Deg
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|23|UN|1|Beam Axial Span
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|24|UN|1|Beam Lateral Min
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|25|UN|1|Beam Lateral Span
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|26|UN|1|Beam Axial Min
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|27|UN|1|Num Display Samples
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|28|UN|1|DVolume Width
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|29|UN|1|DVolume Depth
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|30|UN|1|DVolume Height
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|31|UN|1|DVolume Pos X
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|32|UN|1|DVolume Pos Y
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|33|UN|1|DVolume Pos Z
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|34|UN|1|DBeam Axial Min
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|35|UN|1|DBeam Axial Span
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|37|UN|1|DBeam Lateral Span
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|38|UN|1|Number of Volumes in Sequence
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|39|UN|1|DByte Mask Offset
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|40|UN|1|DByte Mask Size
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|50|LO|1|Private Creator Version of Bookmark
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|51|US|1|BCut Plane Enable
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|52|US|1|BMpr Color Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|53|US|1|BMpr Dynamic Range Db
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|54|US|1|BMpr Gray Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|55|US|1|BVolume Render Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|56|US|1|BVr Brightness
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|57|US|1|BVr Contrast
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|58|US|1|BVr Color Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|59|US|1|BVr Dynamic Range Db
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5a|US|1|BVr Gray Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5b|US|1|BVr Gray Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5c|US|1|BVr Threshold High
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5d|US|1|BVr Threshold Low
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5e|US|1|BPre Process Filter Mix
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|5f|US|1|CCut Plane Enable
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|60|US|1|CFront Clip Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|61|US|1|CMpr Color Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|62|US|1|CMpr Color Flow Priority Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|63|US|1|CVolume Render Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|64|US|1|CVr Color Map Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|65|US|1|CVr Color Flow Priority Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|66|US|1|CVr Opacity
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|67|US|1|CVr Threshold High
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|68|US|1|CVr Threshold Low
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|69|US|1|Voi Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6a|US|1|Voi Rotation Offset Deg
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6b|FD|1|Voi Size Ratio X
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6c|FD|1|Voi Size Ratio Y
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6d|FD|1|Voi Size Ratio Z
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6e|US|1|Voi Sync Plane
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|6f|US|1|Voi View Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|70|FD|1-n|Vr Orientation A
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|71|FD|1-n|Mpr Orientation A
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|72|FD|1|Vr Offset Vector
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|73|FD|1|Blending Ratio
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|74|US|1|Fusion Blend Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|75|FD|1|Quality Factor
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|76|US|1|Renderer Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|77|US|1|Slice Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|78|US|1|Active Quad
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|79|US|1|Screen Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7a|US|1|Cut Plane Side
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7b|US|1|Wireframe Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7c|US|1|Crossmark Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7d|US|1|Mpr Display Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7e|US|1|Volume Display Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|7f|US|1|Last Reset
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|80|US|1|Last Non Full Screen Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|81|US|1|Mpr Tool Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|82|US|1|Voi Tool Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|83|US|1|Tool Loop Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|84|US|1|Volume Arb Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|85|US|1|Mpr Zoom Enabled
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|86|US|1|Is Volume Zoom Enabled
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|87|SS|1|Zoom Level Mpr
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|88|SS|1|Zoom Level Volume
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|89|US|1|Is Auto Rotate Enabled
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8a|US|1|Auto Rotate Axis
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8b|US|1|Auto Rotate Range Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8c|US|1|Auto Rotate Speed Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8d|US|1|CVr Brightness
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8e|US|1|CFlow State Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|8f|US|1|BSubmode Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|90|US|1|CSubmode Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|91|US|1|Cut Plane
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|92|US|1|Bookmark Chunk Id
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|93|US|1|Sequence Min Chunk Id
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|94|US|1|Sequence Max Chunk Id
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|95|FD|1|Volume Rate Hz
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9a|FD|1|Voi Position Offset X
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9b|FD|1|Voi Position Offset Y
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9c|FD|1|Voi Position Offset Z
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9d|US|1|Vr Tool Index
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9e|US|1|Shading Percent
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|9f|US|1|Volume Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|a0|US|1|Vr Quad Display Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|a1|FD|1-n|Mpr Center Location
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e0|US|1|Slice Range Type
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e1|US|1|Slice MPR Plane
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e2|US|1|Slice Layout
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e3|FD|1|Slice Spacing
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e4|US|1|Thin Vr Mode
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e5|US|1|Thin Vr Thickness
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e6|FD|1|Curved TOP VOI Pivot X
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e7|FD|1|Curved TOP VOI Pivot Y
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e8|FD|1|Curved TOP VOI Pivot Z
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|e9|US|1|Curved TOP VOI Quadrant
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|ea|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|ed|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|ee|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|ef|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f0|US|1-n|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f1|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f2|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f3|US|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f4|FD|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f5|LO|1|Unknown
0039|SIEMENS MED SMS USG ANTARES 3D VOLUME|f6|LT|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|50|LO|1|Private Creator Version of Bookmark
0039|SIEMENS MED SMS USG S2000 3D VOLUME|51|US|1|BCut Plane Enable
0039|SIEMENS MED SMS USG S2000 3D VOLUME|52|US|1|BMpr Color Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|53|US|1|BMpr Dynamic Range Db
0039|SIEMENS MED SMS USG S2000 3D VOLUME|54|US|1|BMpr Gray Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|55|US|1|BVolume Render Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|56|US|1|BVr Brightness
0039|SIEMENS MED SMS USG S2000 3D VOLUME|57|US|1|BVr Contrast
0039|SIEMENS MED SMS USG S2000 3D VOLUME|58|US|1|BVr Color Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|59|US|1|BVr Dynamic Range Db
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5a|US|1|BVr Gray Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5b|US|1|BVr Gray Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5c|US|1|BVr Threshold High
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5d|US|1|BVr Threshold Low
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5e|US|1|BPre Process Filter Mix
0039|SIEMENS MED SMS USG S2000 3D VOLUME|5f|US|1|CCut Plane Enable
0039|SIEMENS MED SMS USG S2000 3D VOLUME|60|US|1|CFront Clip Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|61|US|1|CMpr Color Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|62|US|1|CMpr Color Flow Priority Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|63|US|1|CVolume Render Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|64|US|1|CVr Color Map Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|65|US|1|CVr Color Flow Priority Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|66|US|1|CVr Opacity
0039|SIEMENS MED SMS USG S2000 3D VOLUME|67|US|1|CVr Threshold High
0039|SIEMENS MED SMS USG S2000 3D VOLUME|68|US|1|CVr Threshold Low
0039|SIEMENS MED SMS USG S2000 3D VOLUME|69|US|1|Voi Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6a|US|1|Voi Rotation Offset Deg
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6b|FD|1|Voi Size Ratio X
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6c|FD|1|Voi Size Ratio Y
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6d|FD|1|Voi Size Ratio Z
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6e|US|1|Voi Sync Plane
0039|SIEMENS MED SMS USG S2000 3D VOLUME|6f|US|1|Voi View Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|70|FD|1-n|Vr Orientation A
0039|SIEMENS MED SMS USG S2000 3D VOLUME|71|FD|1-n|Mpr Orientation A
0039|SIEMENS MED SMS USG S2000 3D VOLUME|72|FD|1|Vr Offset Vector
0039|SIEMENS MED SMS USG S2000 3D VOLUME|73|FD|1|Blending Ratio
0039|SIEMENS MED SMS USG S2000 3D VOLUME|74|US|1|Fusion Blend Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|75|FD|1|Quality Factor
0039|SIEMENS MED SMS USG S2000 3D VOLUME|76|US|1|Renderer Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|77|US|1|Slice Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|78|US|1|Active Quad
0039|SIEMENS MED SMS USG S2000 3D VOLUME|79|US|1|Screen Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7a|US|1|Cut Plane Side
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7b|US|1|Wireframe Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7c|US|1|Crossmark Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7d|US|1|Mpr Display Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7e|US|1|Volume Display Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|7f|US|1|Last Reset
0039|SIEMENS MED SMS USG S2000 3D VOLUME|80|US|1|Last Non Full Screen Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|81|US|1|Mpr Tool Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|82|US|1|Voi Tool Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|83|US|1|Tool Loop Mode
0119|MRSC|1225|DS|1-n|PercentileLimits
0039|SIEMENS MED SMS USG S2000 3D VOLUME|84|US|1|Volume Arb Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|85|US|1|Mpr Zoom Enabled
0039|SIEMENS MED SMS USG S2000 3D VOLUME|86|US|1|Is Volume Zoom Enabled
0039|SIEMENS MED SMS USG S2000 3D VOLUME|87|SS|1|Zoom Level Mpr
0039|SIEMENS MED SMS USG S2000 3D VOLUME|88|SS|1|Zoom Level Volume
0039|SIEMENS MED SMS USG S2000 3D VOLUME|89|US|1|Is Auto Rotate Enabled
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8a|US|1|Auto Rotate Axis
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8b|US|1|Auto Rotate Range Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8c|US|1|Auto Rotate Speed Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8d|US|1|CVr Brightness
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8e|US|1|CFlow State Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|8f|US|1|BSubmode Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|90|US|1|CSubmode Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|91|US|1|Cut Plane
0039|SIEMENS MED SMS USG S2000 3D VOLUME|92|US|1|Bookmark Chunk Id
0039|SIEMENS MED SMS USG S2000 3D VOLUME|93|US|1|Sequence Min Chunk Id
0039|SIEMENS MED SMS USG S2000 3D VOLUME|94|US|1|Sequence Max Chunk Id
0039|SIEMENS MED SMS USG S2000 3D VOLUME|95|FD|1|Volume Rate Hz
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9a|FD|1|Voi Position Offset X
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9b|FD|1|Voi Position Offset Y
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9c|FD|1|Voi Position Offset Z
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9d|US|1|Vr Tool Index
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9e|US|1|Shading Percent
0039|SIEMENS MED SMS USG S2000 3D VOLUME|9f|US|1|Volume Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|a0|US|1|Vr Quad Display Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|a1|FD|1-n|Mpr Center Location
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e0|US|1|Slice Range Type
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e1|US|1|Slice MPR Plane
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e2|US|1|Slice Layout
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e3|FD|1|Slice Spacing
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e4|US|1|Thin Vr Mode
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e5|US|1|Thin Vr Thickness
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e6|FD|1|Curved TOP VOI Pivot X
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e7|FD|1|Curved TOP VOI Pivot Y
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e8|FD|1|Curved TOP VOI Pivot Z
0039|SIEMENS MED SMS USG S2000 3D VOLUME|e9|US|1|Curved TOP VOI Quadrant
0039|SIEMENS MED SMS USG S2000 3D VOLUME|ea|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|ed|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|ee|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|ef|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f0|US|1-n|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f1|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f2|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f3|US|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f4|FD|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f5|LO|1|Unknown
0039|SIEMENS MED SMS USG S2000 3D VOLUME|f6|LT|1|Unknown
0039|SIEMENS MED OCS BEAM DISPLAY INFO|76|CS|1|Beam Display Properties
0039|SIEMENS MED OCS PUBLIC RT PLAN ATTRIBUTES|01|UT|1|External Attributes
0039|SIEMENS MED OCS SS VERSION INFO|76|LO|1|Structure Set Predecessor
0011|BioPri3D|20|UL|1|Unknown
0011|BioPri3D|24|DS|1-n|Unknown
0011|BioPri3D|30|LO|1|Unknown
0011|BioPri3D|31|UL|1|Unknown
0011|BioPri3D|32|SL|1|Unknown
0011|BioPri3D|39|CS|1|Unknown
0011|BioPri3D|3a|UL|1|Unknown
0011|BioPri3D|d0|OB|1|Unknown
0011|BioPri3D|e0|UL|1|Unknown
0011|BioPri3D|e1|UL|1|Unknown
0011|BioPri3D|e2|UL|1|Unknown
0011|BioPri3D|e3|US|1|Unknown
0011|BioPri3D|e4|US|1|Unknown
0011|BioPri3D|e5|CS|1|Unknown
0063|BioPri3D|0c|DS|1-n|Unknown
0063|BioPri3D|35|SQ|1|Unknown
0063|BioPri3D|20|US|1|Unknown
0063|BioPri3D|21|UL|1|Unknown
2121|PMI Private Calibration Module Version 2.0|01|ST|1|Calibration Method
2121|PMI Private Calibration Module Version 2.0|02|ST|1|Calibration Method Info
2121|PMI Private Calibration Module Version 2.0|03|FL|1|Calibration Object Size
2121|PMI Private Calibration Module Version 2.0|04|FL|1|Calibration Object S Dev
2121|PMI Private Calibration Module Version 2.0|05|FL|1|Calibration Horizontal Pixel Spacing
2121|PMI Private Calibration Module Version 2.0|06|FL|1|Calibration Vertical Pixel Spacing
2121|PMI Private Calibration Module Version 2.0|08|ST|1|Calibration File Name
2121|PMI Private Calibration Module Version 2.0|09|IS|1|Calibration Frame Number
2121|PMI Private Calibration Module Version 2.0|0a|SH|1|Calibration Object Unit
2121|PMI Private Calibration Module Version 2.0|0b|SS|1|Averaged Calibrations Performed
2121|PMI Private Calibration Module Version 2.0|0c|FL|1|Auto Magnify Factor
2121|PMI Private Calibration Module Version 2.0|0d|FL|1|Horizontal Pixel S Dev
2121|PMI Private Calibration Module Version 2.0|0e|FL|1|Vertical Pixel S Dev
0029|CARDIO-D.R. 1.0|ac|FL|1|Displayed Area Bottom Right Hand Corner Fractional
0029|CARDIO-D.R. 1.0|ad|FL|1|Displayed Area Top Left Hand Corner Fractional
0009|POLYTRON-SMS 2.5|02|OB|1|Unknown
0009|POLYTRON-SMS 2.5|04|OB|1|Unknown
0009|POLYTRON-SMS 2.5|06|OB|1|Unknown
0089|POLYTRON-SMS 2.5|10|OB|1|Unknown
300b|SIEMENS MED SYNGO RT|10|CS|1|Plan Type
300b|SIEMENS MED SYNGO RT|11|LT|1|Delivery Warning Dose Comment
300b|SIEMENS MED SYNGO RT|12|LO|1|Imager Organ Program
300b|SIEMENS MED SYNGO RT|13|DS|1|XA Image SID
300b|SIEMENS MED SYNGO RT|14|DS|1|XA Image Receptor Angle
300b|SIEMENS MED SYNGO RT|15|CS|1|Target Prescription Dose Type
300b|SIEMENS MED SYNGO RT|16|IS|1|Referenced Target ROI Number
300b|SIEMENS MED SYNGO RT|17|UT|1|RT Private Data
300b|SIEMENS MED SYNGO RT|18|SQ|1|Referenced Siemens Non Image Sequence
300b|SIEMENS MED SYNGO RT|19|CS|1|Verification Method
300b|SIEMENS MED SYNGO RT|20|SQ|1|Alternative Treatment Machine Name Sequence
300b|SIEMENS MED SYNGO RT|24|DS|1|Imager Angular Angle
300b|SIEMENS MED SYNGO RT|25|DS|1|Imager Isocentric Angle
300b|SIEMENS MED SYNGO RT|26|DS|1|Imager Vertical Position
300b|SIEMENS MED SYNGO RT|27|DS|1|Imager Longitudinal Position
300b|SIEMENS MED SYNGO RT|28|DS|1|Imager Lateral Position
300b|SIEMENS MED SYNGO RT|29|CS|1|Imager Angular Rotation Direction
300b|SIEMENS MED SYNGO RT|2a|CS|1|Imager Isocentric Rotation Direction
300b|SIEMENS MED SYNGO RT|2b|DS|1|Requested Scanning Spot Size
300b|SIEMENS MED SYNGO RT|2c|DS|1|Imager Orbital Angle
300b|SIEMENS MED SYNGO RT|2e|CS|1|Imaging Technique
300b|SIEMENS MED SYNGO RT|2f|CS|1|Imager Orbital Rotation Direction
300b|SIEMENS MED SYNGO RT|30|LO|1|Patient Barcode
300b|SIEMENS MED SYNGO RT|31|SH|3|Beam Modifier Type
300b|SIEMENS MED SYNGO RT|32|FL|3|Source to Range Shifter Distance
300b|SIEMENS MED SYNGO RT|33|SH|3|Treatment Room Name
300b|SIEMENS MED SYNGO RT|60|IS|1-n|Ordered Referenced Beam Numbers
300b|SIEMENS MED SYNGO RT|66|LT|1|Fraction Delivery Notes
300b|SIEMENS MED SYNGO RT|67|LO|1|Record ID
300b|SIEMENS MED SYNGO RT|76|CS|1|Fraction Group Code
300b|SIEMENS MED SYNGO RT|77|IS|1|Referenced Treatment Beam Number
300b|SIEMENS MED SYNGO RT|78|DS|1|Fraction Dose to Dose Reference
300b|SIEMENS MED SYNGO RT|80|SQ|1|Referenced Target ROI Sequence
300b|SIEMENS MED SYNGO RT|82|DS|1|Target ROI Lateral Expansion Margin
300b|SIEMENS MED SYNGO RT|83|DS|1|Target ROI Distal Expansion Margin
300b|SIEMENS MED SYNGO RT|84|DS|1|Target ROI Proximal Expansion Margin
300b|SIEMENS MED SYNGO RT|85|DS|2|Scan Grid Lateral Distance
300b|SIEMENS MED SYNGO RT|86|DS|1|Scan Grid Longitudinal Distance
300b|SIEMENS MED SYNGO RT|87|DS|1|Beam Weight
300b|SIEMENS MED SYNGO RT|89|DS|3|Point on Plane
300b|SIEMENS MED SYNGO RT|8a|DS|3|Norm Vector of Plane
300b|SIEMENS MED SYNGO RT|8b|DS|1|Plane Thickness
300b|SIEMENS MED SYNGO RT|90|SQ|1|Treatment Approval Sequence
300b|SIEMENS MED SYNGO RT|98|DS|1|Treatment Room Temperature
300b|SIEMENS MED SYNGO RT|99|DS|1|Treatment Room Air Pressure
300b|SIEMENS MED SYNGO RT|9b|SQ|1|Split Plane Sequence
300b|SIEMENS MED SYNGO RT|9c|IS|1|Display Color
300b|SIEMENS MED SYNGO RT|9d|SH|1|Beam Group Name
300b|SIEMENS MED SYNGO RT|a0|DT|1|Expire DateTime
300b|SIEMENS MED SYNGO RT|a1|OB|1|Checksum Encryption Code
300b|SIEMENS MED SYNGO RT|a2|CS|1|Setup Type
300b|SIEMENS MED SYNGO RT|a3|IS|1|Number of Therapy Detectors
300b|SIEMENS MED SYNGO RT|a4|SQ|1|Therapy Detector Sequence
300b|SIEMENS MED SYNGO RT|a5|IS|1|Therapy Detector Number
300b|SIEMENS MED SYNGO RT|a6|SH|1|Therapy Detector Setup ID
300b|SIEMENS MED SYNGO RT|a7|SQ|1|Therapy Detector Settings Sequence
300b|SIEMENS MED SYNGO RT|a8|IS|1|Referenced Therapy Detector Number
300b|SIEMENS MED SYNGO RT|a9|DS|1|Therapy Detector Position
300b|SIEMENS MED SYNGO RT|b0|IS|1|Scan Spot Resumption Index
300b|SIEMENS MED SYNGO RT|b1|OW|1|Phantom Detector Measurements
300b|SIEMENS MED SYNGO RT|b2|UT|1|Treatment Events
300b|SIEMENS MED SYNGO RT|c0|SQ|1|Dose Optimization Constraint Sequence
300b|SIEMENS MED SYNGO RT|c8|DS|1|Target Maximum Dose Constraint
300b|SIEMENS MED SYNGO RT|c9|DS|1|Target Maximum Dose Constraint Weight
300b|SIEMENS MED SYNGO RT|ca|DS|1|Target Minimum Dose Constraint
300b|SIEMENS MED SYNGO RT|cb|DS|1|Target Minimum Dose Constraint Weight
300b|SIEMENS MED SYNGO RT|cc|DS|1|Organ At Risk Maximum Dose Constraint
300b|SIEMENS MED SYNGO RT|cd|DS|1|Organ At Risk Maximum Dose Constraint Weight
300b|SIEMENS MED SYNGO RT|ce|SQ|1|DVH Constraint Sequence
300b|SIEMENS MED SYNGO RT|cf|DS|1|DVH Constraint Volume Limit
300b|SIEMENS MED SYNGO RT|d0|CS|1|DVH Constraint Volume Units
300b|SIEMENS MED SYNGO RT|d1|DS|1|DVH Constraint Dose Limit
300b|SIEMENS MED SYNGO RT|d3|CS|1|DVH Constraint Direction
300b|SIEMENS MED SYNGO RT|d4|DS|1|DVH Constraint Weight
300b|SIEMENS MED SYNGO RT|d5|CS|1|Optimized Dose Type
300b|SIEMENS MED SYNGO RT|d6|UT|1|Dose Calculation and Optimization Parameters
300b|SIEMENS MED SYNGO RT|d7|DS|1|Applied Renormalization Factor
300b|SIEMENS MED SYNGO RT|d8|CS|1|Dose Constraint Status
300b|SIEMENS MED SYNGO RT|d9|DS|1|Organ At Risk Minimum Dose Constraint
300b|SIEMENS MED SYNGO RT|da|DS|1|Organ At Risk Minimum Dose Constraint Weight
300b|SIEMENS MED SYNGO RT|e0|SQ|1|Base Data Group Sequence
300b|SIEMENS MED SYNGO RT|e1|CS|1|Physics Base Data Group ID
300b|SIEMENS MED SYNGO RT|e2|CS|1|Biological Base Data Group ID
300b|SIEMENS MED SYNGO RT|e3|CS|1|Imaging Base Data Group ID
300b|SIEMENS MED SYNGO RT|e4|CS|1|Dosimetric Base Data Group ID
300b|SIEMENS MED SYNGO RT|e5|OB|1|Configuration Baseline
300b|SIEMENS MED SYNGO RT|e6|OB|1|Configuration Objects
300b|SIEMENS MED SYNGO RT|e7|CS|1|Confidence Measure Units
300b|SIEMENS MED SYNGO RT|e8|DS|1|Confidence Measure Value
300b|SIEMENS MED SYNGO RT|e9|LO|1|Imager Organ Program Name
300b|SIEMENS MED SYNGO RT|eb|CS|1|Body Region
300b|SIEMENS MED SYNGO RT|ec|CS|1|Prefinalized Status
300b|SIEMENS MED SYNGO RT|ed|OB|1|Dosimetric Checksum Encryption Code
300b|SIEMENS MED SYNGO RT|ee|SQ|1|Referenced Report Sequence
300b|SIEMENS MED SYNGO RT|ef|CS|1|Maintain Checksum Compatibility
300b|SIEMENS MED SYNGO RT|f0|DS|1|Dose Statistical Uncertainty
300b|SIEMENS MED SYNGO RT|f1|CS|1|Interpreted Radiation Type
7fd1|SIEMENS SYNGO ULTRA-SOUND TOYON DATA STREAMING|01|OB|1|Padding
7fd1|SIEMENS SYNGO ULTRA-SOUND TOYON DATA STREAMING|09|OB|1|Version ID
7fd1|SIEMENS SYNGO ULTRA-SOUND TOYON DATA STREAMING|10|LO|1|Payload
7fd1|SIEMENS SYNGO ULTRA-SOUND TOYON DATA STREAMING|11|LO|1|After Payload
0021|SIEMENS Ultrasound S2000|00|US|1|Nipple Position
0021|SIEMENS Ultrasound S2000|01|US|1|ABVS Clip Derived From Volume
0079|SMIL_PB79|00|LO|1|Analgesia
0079|SMIL_PB79|01|LO|1|Anesthesia
0079|SMIL_PB79|02|IS|1|Bed Motion
0079|SMIL_PB79|03|LO|1|Food Access
0079|SMIL_PB79|04|DS|1|Histogram Version
0079|SMIL_PB79|06|DS|1|Injection Decay Correction
0079|SMIL_PB79|07|LO|1|Isotope
0079|SMIL_PB79|08|LO|1|Other Drugs
0079|SMIL_PB79|09|IS|1|RebinningType
0079|SMIL_PB79|0a|DS|1|Rebinning Version
0079|SMIL_PB79|0b|IS|1|Reconstruction
0079|SMIL_PB79|0c|DS|1|ReconstructionVersion
0079|SMIL_PB79|0d|LO|1|Injected Compounds
0079|SMIL_PB79|0e|LO|1|Study Model
0079|SMIL_PB79|0f|LO|1|Subject Genus
0079|SMIL_PB79|10|LO|1|Subject Phenotype
0079|SMIL_PB79|11|DS|1|Version
0079|SMIL_PB79|12|LO|1|Water Access
0079|SMIL_PB79|13|DS|1|X Offset
0079|SMIL_PB79|14|DS|1|Y Offset
0079|SMIL_PB79|15|DS|1|Zoom
0079|SMIL_PB79|17|IS|1|Subject Orientation
007b|SMIO_PB7B|00|LO|1|Units
007d|SMIO_PB7D|01|UL|1|Geometry
007d|SMIO_PB7D|02|FL|1|Spacing
007d|SMIO_PB7D|03|FL|1|Origin
0009|TOSHIBA_MEC_OT3|00|LO|1|HIS/RIS Study ID
0029|TOSHIBA MDW NON-IMAGE|08|CS|1|Non-Image Header Type
0029|TOSHIBA MDW NON-IMAGE|09|LO|1|Non-Image Header Version
0029|TOSHIBA MDW NON-IMAGE|20|OB|1|Unknown
0029|TOSHIBA MDW HEADER|08|CS|1|Image Header Type
0029|TOSHIBA MDW HEADER|09|LO|1|Image Header Version
0029|TOSHIBA MDW HEADER|10|OB|1|Image Header Info
0029|TOSHIBA MDW HEADER|18|CS|1|Series Header Type
0029|TOSHIBA MDW HEADER|19|LO|1|Series Header Version
0029|TOSHIBA MDW HEADER|20|OB|1|Series Header Info
0029|TOSHIBA COMAPL HEADER|08|CS|1|COMAPL Header Type
0029|TOSHIBA COMAPL HEADER|09|LO|1|COMAPL Header Version
0029|TOSHIBA COMAPL HEADER|10|OB|1|COMAPL Header Info
0029|TOSHIBA COMAPL HEADER|20|OB|1|COMAPL History Information
0029|TOSHIBA COMAPL HEADER|31|LO|1|Unknown
0029|TOSHIBA COMAPL HEADER|34|LO|1|Unknown
0029|TOSHIBA COMAPL OOG|08|CS|1|COMAPL OOG Type
0029|TOSHIBA COMAPL OOG|09|LO|1|COMAPL OOG Version
0009|MMCPrivate|1c|OB|1|ProtocolAppData
0029|TOSHIBA COMAPL OOG|10|OB|1|COMAPL OOG Info
0029|PMTF INFORMATION DATA|01|SQ|1|Unknown
0029|PMTF INFORMATION DATA|31|LO|1|PMTF Information 1
0029|PMTF INFORMATION DATA|32|UL|1|PMTF Information 2
0029|PMTF INFORMATION DATA|33|UL|1|PMTF Information 3
0029|PMTF INFORMATION DATA|34|CS|1|PMTF Information 4
0029|PMTF INFORMATION DATA|89|LO|1|Unknown
0029|PMTF INFORMATION DATA|90|OB|1|Unknown
7005|TOSHIBA_MEC_CT3|61|LO|1|Synchronized Signal Information
7005|TOSHIBA_MEC_CT3|62|DS|1|Total Raw Data Size
7005|TOSHIBA_MEC_CT3|63|FD|1|CTDIw
7005|TOSHIBA_MEC_CT3|67|UI|1|Volume UID of 4D-Volume
7005|TOSHIBA_MEC_CT3|68|US|1|Total Frame Count in 4D-Volume
7005|TOSHIBA_MEC_CT3|69|US|1|Frame Number in 4D-Volume
7005|TOSHIBA_MEC_CT3|6a|DS|3|Image Position of 4D-Volume Top
7005|TOSHIBA_MEC_CT3|6b|DS|3|Image Position of 4D-Volume Top (Equipment)
7005|TOSHIBA_MEC_CT3|6c|UI|1|SOP Instance UID of 4D-Volume
7005|TOSHIBA_MEC_CT3|6d|UI|1|Series Instance UID of 4D-Volume
7015|TOSHIBA ENCRYPTED SR DATA|00|OB|1|Unknown
7015|TOSHIBA_SR|10|OB|1|Unknown
7015|TOSHIBA_SR|60|OB|1|Unknown
7015|PMTF INFORMATION DATA|73|SQ|1|Unknown
7079|TOSHIBA_MEC_XA3|21|SH|5|Unknown
7079|TOSHIBA_MEC_XA3|22|IS|2|Unknown
7079|TOSHIBA_MEC_XA3|23|IS|2|Unknown
7079|TOSHIBA_MEC_XA3|24|DS|1|Unknown
7079|TOSHIBA_MEC_XA3|25|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|26|DS|2|Unknown
7079|TOSHIBA_MEC_XA3|27|US|2|Unknown
7079|TOSHIBA_MEC_XA3|28|US|1|Unknown
7079|TOSHIBA_MEC_XA3|2a|US|5|Unknown
7079|TOSHIBA_MEC_XA3|2c|SH|3|Unknown
7079|TOSHIBA_MEC_XA3|2d|SS|2|Unknown
7079|TOSHIBA_MEC_XA3|2e|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|2f|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|30|US|1|Unknown
7079|TOSHIBA_MEC_XA3|31|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|32|SH|2|Unknown
7079|TOSHIBA_MEC_XA3|33|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|34|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|35|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|36|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|37|US|4|Unknown
7079|TOSHIBA_MEC_XA3|38|SS|1-n|Unknown
7079|TOSHIBA_MEC_XA3|39|SS|1-n|Unknown
7079|TOSHIBA_MEC_XA3|3a|US|2|Unknown
7079|TOSHIBA_MEC_XA3|3b|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|3c|DS|2|Unknown
7079|TOSHIBA_MEC_XA3|3d|SS|2|Unknown
7079|TOSHIBA_MEC_XA3|3e|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|3f|US|2|Unknown
7079|TOSHIBA_MEC_XA3|40|SH|2|Unknown
7079|TOSHIBA_MEC_XA3|41|SS|2|Unknown
7079|TOSHIBA_MEC_XA3|42|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|43|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|44|US|1|Unknown
7079|TOSHIBA_MEC_XA3|45|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|46|SS|1|Unknown
7079|TOSHIBA_MEC_XA3|47|SS|18|Unknown
7079|TOSHIBA_MEC_XA3|48|US|12|Unknown
7079|TOSHIBA_MEC_XA3|49|US|3|Unknown
7079|TOSHIBA_MEC_XA3|4a|US|1|Unknown
7079|TOSHIBA_MEC_XA3|4b|LO|3|Unknown
7079|TOSHIBA_MEC_XA3|4c|OB|1|Unknown
7079|TOSHIBA_MEC_XA3|4d|SH|3|Unknown
7079|TOSHIBA_MEC_XA3|4e|SL|35|Unknown
7079|TOSHIBA_MEC_XA3|4f|SH|3|Unknown
7079|TOSHIBA_MEC_XA3|50|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|51|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|52|US|1|Unknown
7079|TOSHIBA_MEC_XA3|53|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|54|US|5|Unknown
7079|TOSHIBA_MEC_XA3|55|UL|47-47n|Unknown
7079|TOSHIBA_MEC_XA3|56|US|1|Unknown
7079|TOSHIBA_MEC_XA3|57|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|58|US|1|Unknown
7079|TOSHIBA_MEC_XA3|59|US|2-2n|Unknown
7079|TOSHIBA_MEC_XA3|5a|US|1|Unknown
7079|TOSHIBA_MEC_XA3|5b|US|2|Unknown
7079|TOSHIBA_MEC_XA3|5c|US|2-2n|Unknown
7079|TOSHIBA_MEC_XA3|5d|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|5e|US|2|Unknown
7079|TOSHIBA_MEC_XA3|5f|SS|4-4n|Unknown
7079|TOSHIBA_MEC_XA3|60|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|61|SS|30-30n|Unknown
7079|TOSHIBA_MEC_XA3|62|US|4|Unknown
7079|TOSHIBA_MEC_XA3|63|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|64|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|65|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|66|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|67|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|68|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|69|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|6a|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|6b|US|1-n|Unknown
7079|TOSHIBA_MEC_XA3|6c|US|1|Unknown
7079|TOSHIBA_MEC_XA3|6d|DS|1|Unknown
7079|TOSHIBA_MEC_XA3|6e|LO|1|Unknown
7079|TOSHIBA_MEC_XA3|6f|DS|1|Unknown
7079|TOSHIBA_MEC_XA3|70|DS|1|Unknown
7079|TOSHIBA_MEC_XA3|71|DS|1-n|Unknown
7079|TOSHIBA_MEC_XA3|72|DS|1-n|Unknown
7079|TOSHIBA_MEC_XA3|73|SL|4|Unknown
7079|TOSHIBA_MEC_XA3|74|SL|28|Unknown
7079|TOSHIBA_MEC_XA3|75|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|76|US|1|Unknown
7079|TOSHIBA_MEC_XA3|77|SL|1|Unknown
7079|TOSHIBA_MEC_XA3|78|US|1|Unknown
7079|TOSHIBA_MEC_XA3|79|US|1|Unknown
7079|TOSHIBA_MEC_XA3|7b|SH|1|Unknown
7079|TOSHIBA_MEC_XA3|80|LO|1|Unknown
0009|FDMS 1.0|04|SH|1|ImageControlUnit
0009|FDMS 1.0|06|OW|1|RouteImage UID
0009|FDMS 1.0|0c|OW|1|Film UID
0009|FDMS 1.0|f0|CS|1|Blackening Process Flag
0009|GEMS_IDEN_01|01|LO|1|FullFidelity
0009|GEMS_PETD_01|01|LO|2|Implementation Version Name
0009|GEMS_PETD_01|0b|SH|1|Scan Compatible Version
0009|GEMS_PETD_01|21|SL|1|Count Rate Period
0009|GEMS_PETD_01|29|FL|1|Gantry Tilt Angle
0009|GEMS_PETD_01|3c|FL|1|Post Injected Activity
0009|GEMS_PETD_01|51|SL|1|Upper Coinc Limit
0009|GEMS_PETD_01|5e|UI|1|exam_id
0009|GEMS_PETD_01|60|SH|1|compatible_version
0009|GEMS_PETD_01|79|SH|1|Image Set Compatible Version
0009|GEMS_PETD_01|94|SL|1|Atten Smooth Param
0009|GEMS_PETD_01|9b|FL|1|CAC Skull Offset
0009|GEMS_PETD_01|9f|SL|1|Axial Filter 3D
0009|GEMS_PETD_01|b6|SS|1|IR Loop Filter
0009|GEMS_PETD_01|cd|FL|1|vqc_y_axis_trans
0009|GEMS_PETD_01|da|ST|1|where_is_list_frame
0009|GEMS_PETD_01|db|SL|1|ir_z_filter_flag
0009|GEMS_PETD_01|f0|UI|1|Reformat group
0009|GEMS_PETD_01|f1|SL|1|PET prompt gamma
0009|GEMS_PETD_01|f2|UI|1|PET tracerInjection_UID
0009|GE_YMS_NJ001|31|SH|1|Mobile Location Code
0009|MMCPrivate|01|LO|1|Technologist
0009|MMCPrivate|04|UI|1|ProtocolObjectID
0009|MMCPrivate|05|LO|1|Name
0009|MMCPrivate|06|IS|1|Frequency
0009|MMCPrivate|07|SH|1|UpdateFlag
0009|MMCPrivate|08|SH|1|Directory
0009|MMCPrivate|09|LO|1|Comments
0009|MMCPrivate|0a|LO|1|Region
0009|MMCPrivate|0b|SH|1|Laterality
0009|MMCPrivate|0c|TM|1|TotalScanTime
0009|MMCPrivate|0d|LO|1|ContrastMedium
0009|MMCPrivate|0e|LO|1|CreateDateTime
0009|MMCPrivate|0f|LO|1|Creator
0009|MMCPrivate|10|LO|1|SiteName
0009|MMCPrivate|11|LO|1|ReferringPhysician
0009|MMCPrivate|12|LO|1|Radiologist
0009|MMCPrivate|13|LO|1|Technologist
0009|MMCPrivate|14|UI|1|ProtocolUid
0009|MMCPrivate|15|SH|1|IsInLibrary
0009|MMCPrivate|16|LO|1|Gating
0009|MMCPrivate|17|ST|1|Note
0009|MMCPrivate|18|IS|1|NumberOfTasks
0009|MMCPrivate|19|SH|1|IsFlagRaised
0009|MMCPrivate|1a|SH|1|IsArchived
0009|MMCPrivate|1b|SH|1|IsDefault
0009|MMCPrivate|20|UI|1|TaskInfoObjectID
0009|MMCPrivate|21|LO|1|Name
0009|MMCPrivate|22|SH|1|TaskStatus
0009|MMCPrivate|23|SH|1|TaskPriority
0009|MMCPrivate|24|SH|1|Leaf
0009|MMCPrivate|25|LO|1|TaskID
0009|MMCPrivate|26|IS|1|Frequency
0009|MMCPrivate|27|SH|1|UpdateFlag
0009|MMCPrivate|28|SH|1|Directory
0009|MMCPrivate|29|LO|1|Comments
0009|MMCPrivate|2a|SH|1|Category
0009|MMCPrivate|2b|LO|1|Region
0009|MMCPrivate|2c|SH|1|Laterality
0009|MMCPrivate|2d|TM|1|ScanTime
0009|MMCPrivate|2e|LO|1|ContrastMedium
0009|MMCPrivate|2f|LO|1|CreateDateTime
0009|MMCPrivate|30|LO|1|Creator
0009|MMCPrivate|31|LO|1|SiteName
0009|MMCPrivate|32|LO|1|ReferringPhysician
0009|MMCPrivate|33|LO|1|Radiologist
0009|MMCPrivate|34|LO|1|Technologist
0009|MMCPrivate|35|UI|1|TaskUid
0009|MMCPrivate|36|UI|1|TaskInfoUid
0009|MMCPrivate|37|SH|1|IsInLibrary
0009|MMCPrivate|38|IS|1|TaskOrder
0009|MMCPrivate|39|LO|1|Gating
0009|MMCPrivate|3a|SH|1|Plane
0009|MMCPrivate|3b|LO|1|SequenceType
0009|MMCPrivate|3c|SH|1|IsExecutive
0009|MMCPrivate|3d|ST|1|Note
0009|MMCPrivate|3e|SH|1|AutoStart
0009|MMCPrivate|3f|SH|1|AutoSave
0009|MMCPrivate|40|SH|1|AutoArchive
0009|MMCPrivate|41|IS|1|QueueGroupID
0009|MMCPrivate|42|SH|1|IsFlagRaised
0009|MMCPrivate|43|SH|1|IsArchived
0009|MMCPrivate|44|SH|1|IsDefault
0009|MMCPrivate|45|OB|1|TaskInfoAppData
0009|MMCPrivate|46|SH|1|IsAllowCascadeSave
0009|MMCPrivate|47|SH|1|IsAllowCascadeProtect
0009|MMCPrivate|5f|UI|1|ProtocolObjectID
0009|MMCPrivate|60|OB|1|TaskInfoAppData
0009|MMCPrivate|72|UI|1|ProtocolTaskInfoObjectID
0009|MMCPrivate|73|IS|1|ProtocolTaskOrder
0009|MMCPrivate|74|UI|1|ProtocolTaskUid
0009|MMCPrivate|75|OB|1|ProtocolTaskAppData
0009|MMCPrivate|76|SH|1|ProtocolTaskIsAllowCascadeSave
0009|MMCPrivate|77|SH|1|ProtocolTaskIsAllowCascadeProtect
0011|GEMS_PATI_01|10|SS|1|PatientStatus
0011|GEMS_PETD_01|02|UI|1|PET ROI.roi_id
0011|GEMS_PETD_01|03|UI|1|PET ROI.image_id
0011|GEMS_PETD_01|04|UI|1|PET ROI.compatible_version
0011|GEMS_PETD_01|05|SH|1|PET ROI.software_version
0011|GEMS_PETD_01|06|LO|1|PET ROI.roi_name
0011|GEMS_PETD_01|07|DT|1|PET ROI.roi_datetime
0011|GEMS_PETD_01|08|SL|1|PET ROI.roi_type
0011|GEMS_PETD_01|09|FL|1|PET ROI.center_x
0011|GEMS_PETD_01|0a|FL|1|PET ROI.center_y
0011|GEMS_PETD_01|0b|FL|1|PET ROI.width
0011|GEMS_PETD_01|0c|FL|1|PET ROI.height
0011|GEMS_PETD_01|0d|FL|1|PET ROI.angle
0011|GEMS_PETD_01|0e|SL|1|PET ROI.number_of_points
0011|GEMS_PETD_01|0f|OB|1|PET ROI.roi_data
0011|GEMS_PETD_01|10|SL|1|PET ROI.roi_size
0011|GEMS_PETD_01|11|LO|1|PET ROI.color
0011|GEMS_PETD_01|12|SL|1|PET ROI.line_type
0011|GEMS_PETD_01|13|SL|1|PET ROI.line_width
0011|GEMS_PETD_01|14|SL|1|PET ROI.roi_number
0011|GEMS_PETD_01|15|SL|1|PET ROI.convex
0011|GEMS_PETD_01|16|SL|1|PET ROI.atten_cor_flag
0013|CTP|10|LO|1|Project Name
0013|CTP|14|UN|1|Visibility
0013|GEMS_PETD_01|02|UI|1|PET Annotation.annotation_id
0013|GEMS_PETD_01|03|UI|1|PET Annotation.image_id
0013|GEMS_PETD_01|04|SH|1|PET Annotation.compatible_version
0013|GEMS_PETD_01|05|SH|1|PET Annotation.software_version
0013|GEMS_PETD_01|06|SL|1|PET Annotation.type
0013|GEMS_PETD_01|07|LO|1|PET Annotation.font_name
0013|GEMS_PETD_01|08|SH|1|PET Annotation.font_size
0013|GEMS_PETD_01|09|LO|1|PET Annotation.foreground_color
0013|GEMS_PETD_01|0a|LO|1|PET Annotation.background_color
0013|GEMS_PETD_01|0b|SL|1|PET Annotation.coordinate_system
0013|GEMS_PETD_01|0c|FL|1|PET Annotation.start_x
0013|GEMS_PETD_01|0d|FL|1|PET Annotation.start_y
0013|GEMS_PETD_01|0e|FL|1|PET Annotation.end_x
0013|GEMS_PETD_01|0f|FL|1|PET Annotation.end_y
0013|GEMS_PETD_01|10|SL|1|PET Annotation.start_symbol
0013|GEMS_PETD_01|11|SL|1|PET Annotation.end_symbol
0013|GEMS_PETD_01|12|OB|1|PET Annotation.annotation_data
0013|GEMS_PETD_01|13|SL|1|PET Annotation.annotation.size
0013|GEMS_PETD_01|14|LO|1|PET Annotation.label_id
0015|GEMS_PETD_01|1a|US|1|Physio Gating Type
0015|GEMS_PETD_01|1b|US|1|Total Number of Bins
0015|GEMS_PETD_01|1c|US|1|% Phase Value
0015|GEMS_PETD_01|1d|SL|1|Phase Matched Series
0015|GEMS_PETD_01|1e|SL|1|CTAC Percent Value
0015|GEMS_PETD_01|1f|UL|1|PET Recon Parameters Exists
0015|GEMS_PETD_01|20|SL|1|First Packet Number
0015|GEMS_PETD_01|21|FL|1|IR Loop Filter Ratio
0015|GEMS_PETD_01|22|FL|1|IR Loop Filter Correction
0015|GEMS_PETD_01|23|UL|1|BP3d Filter FlagU
0015|GEMS_PETD_01|24|FL|1|BP3d Filter CutoffU
0015|GEMS_PETD_01|25|SL|1|BP3d Filter OrderU
0015|GEMS_PETD_01|26|UL|1|BP3d Filter FlagV
0015|GEMS_PETD_01|27|FL|1|BP3d Filter OrderV
0015|GEMS_PETD_01|28|SL|1|BP3d Filter CutoffV
0015|GEMS_PETD_01|29|UL|1|Decay Flag
0015|GEMS_PETD_01|2e|UL|1|Image filter 3d flag
0015|GEMS_PETD_01|2f|UL|1|WCC Cal Flag
0015|GEMS_PETD_01|30|UL|1|Emission Scatter Flag
0015|GEMS_PETD_01|31|UL|1|Recon Algorithm
0015|GEMS_PETD_01|32|UL|1|Normalization Flag
0015|GEMS_PETD_01|33|UL|1|Emission Deadtime Flag
0015|GEMS_PETD_01|34|UL|1|Emission Random Flag
0015|GEMS_PETD_01|35|UL|1|Blank Scan Flag
0119|MRSC|1226|DS|1-n|InPlaneRotation
0015|GEMS_PETD_01|39|SL|1|Event histogram Format
0015|GEMS_PETD_01|3a|SL|1|Number of Detector Rows
0015|GEMS_PETD_01|3b|SL|1|Number of Detector Columns
0015|GEMS_PETD_01|3c|US|1|Recon Matrix Size
0015|GEMS_PETD_01|3d|UL|1|PET Sharp IR Flag
0015|GEMS_PETD_01|3e|UL|1|PET Scatter Limit
0017|GEMS_PETD_01|02|SH|1|compatible_version
0019|ADAC_IMG|02|IS|1|ADAC Pegasys File Size
0019|GEMS_ACQU_01|02|SL|1|NumberOfCellsInDetector
0019|GEMS_ACQU_01|25|SS|1|MidScanFlag
0019|GEMS_ACQU_01|40|SS|1|StatReconFlag
0019|GEMS_ACQU_01|41|SS|1|ComputeType
0019|GEMS_ACQU_01|6a|SS|1|DependantOnNumberOfViewsProcessed
0019|GEMS_ACQU_01|92|SL|1|SliceOffsetOnFrequencyAxis
0019|GEMS_ACQU_01|9e|LO|1|InternalPulseSequenceName
0019|GEMS_ACQU_01|b2|DS|1|UserData
0019|GEMS_ACQU_01|cb|SS|1|PrescribedFlowAxis
0019|GEMS_ACQU_01|dd|SS|1|OverrangeCorrectionUsed
0019|GEMS_PETD_01|09|FL|1|activity_factor_hr
0019|GEMS_PETD_01|18|UI|1|WCC Image Set ID
0019|GE_YMS_NJ001|02|SL|1|Detector Channel
0019|GE_YMS_NJ001|23|DS|1|Table speed
0019|GE_YMS_NJ001|24|DS|1|Mid scan time
0019|GE_YMS_NJ001|26|SL|1|Tube Azimuth
0019|GE_YMS_NJ001|27|DS|1|Gantry Velocity
0019|GE_YMS_NJ001|39|SS|1|SFOV type
0019|GE_YMS_NJ001|42|SS|1|Segment number
0019|GE_YMS_NJ001|43|SS|1|Total segments required
0019|MMCPrivate|04|DS|1|Max Fscalor
0019|MMCPrivate|05|LO|1|Series Category Type
0019|MMCPrivate|09|DS|1|Image Reconstruction Diameter
0019|MMCPrivate|20|UI|1|MultiFrameSopInstanceUid
0019|SIEMENS CT VA0  COAD|90|DS|1|OsteoOffset
0019|SIEMENS CT VA0  COAD|b0|DS|1|Feed per Rotation
0019|SIEMENS CT VA0  COAD|be|DS|1|Expiratoric Reserve Volume
0019|Siemens MED NM|0f|SL|1-n|Siemens ICON Data Type
0019|Siemens MED NM|a5|SS|1-n|Number of repeats per phase
0019|Siemens MED NM|a6|SS|1-n|Cycles per repeat
0019|Siemens MED NM|a7|SL|1-n|Repeat start time
0019|Siemens MED NM|a8|SL|1-n|Repeat stop time
0019|Siemens MED NM|a9|SL|1-n|Effective repeat time
0019|Siemens MED NM|aa|SS|1-n|Acquired cycles per repeat
0021|FDMS 1.0|40|IS|1|ImageNoInTheSet
0021|GEMS_RELA_01|03|SS|1|SeriesFromWhichPrescribed
0021|GEMS_RELA_01|82|DS|1|AutoWindowLevelBeta
0021|GEMS_RELA_01|90|SS|1|TubeFocalSpotPosition
0021|GEMS_RELA_01|92|FL|1|BiopsyTLocation
0021|SIEMENS MED|11|DS|2|Target
0021|Siemens MED NM|00|OB|1|ECAT File Menu Header
0021|Siemens MED NM|01|OB|1|ECAT File Subheader
0023|GEMS_PETD_01|02|0B|1|PET raw_data_blob
0023|GEMS_STDY_01|80|SQ|1|Has MPPS Related Tags
0023|Siemens MED NM|01|US|1|DICOM Reader Flag
0027|GEMS_IMAG_01|1c|SL|1|VmaMamp
0027|GEMS_IMAG_01|44|FL|1|CenterSCoordOfPlaneImage
0119|MRSC|1230|IS|1-n|ReSample
0027|GE_YMS_NJ001|10|SS|1|Scout Type
0027|GE_YMS_NJ001|50|FL|1|Scan start location
0027|GE_YMS_NJ001|51|FL|1|Scan end location
0029|GEMS_CT_FLRO_01|01|SS|1|CT Int Fluoro
0029|GEMS_CT_FLRO_01|02|DS|1|Image Precise Location
0029|GEMS_IMPS_01|06|DS|1|LowerRangeOfPixels
0029|GEMS_IMPS_01|0a|SS|1|LowerRangeOfPixels
0029|MMCPrivate|11|LO|1|Echo Allocation
0029|MMCPrivate|29|DS|1|Table Position
0029|MMCPrivate|2b|DS|1|Navi Final Gate Width
0029|MMCPrivate|2d|DS|1|Navi Final Gate Position
0029|MMCPrivate|48|CS|1|Respiratory Motion Compensation Technique
0029|MMCPrivate|61|LO|1|Window Center and Width Explanation
0029|MMCPrivate|66|CS|1|Inversion Recovery
0029|MMCPrivate|6a|CS|1|Partial Fourier
0029|MMCPrivate|6c|CS|1|ResonantNucleus
0029|MMCPrivate|6d|CS|1|KSpaceFiltering
0029|MMCPrivate|6e|CS|1|ApplicableSafetyStandardAgency
0029|MMCPrivate|6f|LO|1|ApplicableSafetyStandardDescription
0029|MMCPrivate|88|US|1|MRAcquisition Frequency Encoding Steps
0029|MMCPrivate|a2|FD|1|Transmitter Frequency
0029|MMCPrivate|a5|FD|1|Velocity Encoding Direction
0029|MMCPrivate|ab|CS|1|Volumetric Properties
0029|MMCPrivate|c6|DS|1|SelectiveIROrientation
0029|MMCPrivate|c7|LO|1|SelectiveIRThickness
0029|MMCPrivate|c8|SH|1|RephaseOrderSlice
0029|MMCPrivate|c9|SH|1|RephaseOrderPhase
0029|MMCPrivate|ca|SH|1|RephaseOrderFreq
0029|MMCPrivate|cb|ST|1|MetaboliteMapDescription
0029|MMCPrivate|cc|SQ|1|volumeLocalizationSeq
0029|MMCPrivate|cd|FD|1|SlabThickness
0029|MMCPrivate|ce|FD|1|SlabOrientation
0029|MMCPrivate|cf|FD|1|MidSlabPosition
0029|MMCPrivate|d1|LO|1|IRThicknessRatio
0029|MMCPrivate|d2|LO|1|BBIRThicknessRatio
0029|MMCPrivate|d4|IS|1|MultiFrameFrameNumber
0029|SIEMENS CSA ENVELOPE|10|OB|1|syngo Report Data
0029|SIEMENS MEDCOM HEADER|08|CS|1|MedComHeaderType
0029|SIEMENS MEDCOM HEADER|43|LO|1|ApplicationHeaderVersion
0029|SIEMENS MEDCOM HEADER|70|SQ|1|Siemens Link Sequence
0029|SIEMENS MEDCOM HEADER|75|OB|1|Referenced Object Device Location
0033|SIEMENS MED NM|00|FL|1-n|Flood Correction Matrix Detector 1
0033|SIEMENS MED NM|19|FL|1-n|NCO Data for detector 2
0033|SIEMENS MED NM|21|FL|1|Gantry correction angle
0033|SIEMENS MED NM|35|FL|1|Weight Factor Table For Coincidence Acquisitions
0039|GEMS_0039|95|LO|1|Unknown
0040|GEMS_HELIOS_01|19|SS|1|Air Calibration Date
0041|MMCPrivate|01|OB|1|RawDataAppData
0041|MMCPrivate|02|SQ|1|RawDataIndex
0041|MMCPrivate|03|LO|1|ChannelNumber
0041|MMCPrivate|04|LO|1|AxisDirection
0041|MMCPrivate|05|LO|1|SlabNumbe
0041|MMCPrivate|06|LO|1|CardiacPhaseNumbe
0041|MMCPrivate|07|LO|1|EchoNumber
0041|MMCPrivate|08|LO|1|SliceEncodeNumber
0041|MMCPrivate|09|LO|1|NsaNumber
0041|MMCPrivate|0a|OB|1|RawData
0041|MMCPrivate|0b|SS|1|RawDataMRInfo
0041|MMCPrivate|0c|IS|1|NumberOfVoxels
0041|MMCPrivate|0d|DS|1|MixingTime
0041|MMCPrivate|0e|DS|1|ADDiff
0041|MMCPrivate|0f|LO|1|ScanTime
0041|MMCPrivate|10|LO|1|NumPreSat
0041|MMCPrivate|11|LO|1|IsStoredToPortableMedia
0041|MMCPrivate|12|DS|1|Voi1
0041|MMCPrivate|13|DS|1|Voi2
0041|MMCPrivate|14|DS|1|VoxelSize
0041|MMCPrivate|15|IS|1|FreqPoint
0041|MMCPrivate|16|SH|1|LowOrderShim
0041|MMCPrivate|17|SH|1|EccLevel
0041|MMCPrivate|18|FL|1|FwhmHz
0041|MMCPrivate|19|FL|1|FwhmPpm
0041|MMCPrivate|1a|FL|1|WaterSupRate
0043|GEMS_PARM_01|03|SS|1|GradientOffsetInY
0043|GEMS_PARM_01|17|DS|1|IBHImageScaleFactors
0043|GEMS_PARM_01|2d|SH|1|StringSlopField1
0043|GEMS_PARM_01|4e|FL|4|DurationOfXrayOn
0043|GEMS_PARM_01|63|SH|1|Raw Data ID
0043|GEMS_PARM_01|65|US|1|Motion Correction Indicator
0043|GEMS_PARM_01|82|LO|1-n|System Configuration Information
0043|GEMS_PARM_01|8b|OB|1|FMRI Binary Data Block
0043|GEMS_PARM_01|97|LO|8|Image Filtering Parameters
0043|GEMS_PARM_01|9b|DS|1|NPW factor
0043|GEMS_PARM_01|9c|OB|1|Research Tag 1
0043|GEMS_PARM_01|9d|OB|1|Research Tag 2
0043|GEMS_PARM_01|9e|OB|1|Research Tag 3
0043|GEMS_PARM_01|9f|OB|1|Research Tag 4
0043|GEMS_PARM_01|a0|SQ|1|Spectroscopy Pixel Sequence
0043|GEMS_PARM_01|a1|SQ|1|Spectroscopy Default Display Sequence
0043|GEMS_PARM_01|a2|DS|1-n|MEF Data
0043|GEMS_PARM_01|a3|CS|1|ASL Contrast technique
0043|GEMS_PARM_01|a4|LO|1|Detailed text for ASL labeling technique
0043|GEMS_PARM_01|a5|IS|1|Duration of the label or control pulse
0043|GEMS_PARM_01|a6|DS|1|Offset frequency value for FastB1map
0043|GEMS_PARM_01|a7|DS|1|Motion Encoding Factor
0043|GE_YMS_NJ001|12|SS|3|X-Ray Chain
0043|GE_YMS_NJ001|1e|DS|1|Delta start time [msec]
0043|GE_YMS_NJ001|35|US|1|Infant Indicator
0043|GE_YMS_NJ001|37|CS|1|Gantry Type
0043|GE_YMS_NJ001|38|SH|1|Raw data ID
0043|GE_YMS_NJ001|39|IS|1|Reconstruction Matrix
0043|GE_YMS_NJ001|40|CS|1-n|Image Filter
0043|GE_YMS_NJ001|41|US|1|Prospective Addition Indicator
0043|GE_YMS_NJ001|43|US|1|Motion Correction Indicator
0043|GE_YMS_NJ001|44|US|1|Helical Correction Indicator
0043|GE_YMS_NJ001|45|US|1|Cine Correction Indicator
0043|GE_YMS_NJ001|46|US|1|IBO Correction Indicator
0043|GE_YMS_NJ001|47|US|1|BBH Correction Indicator
0043|GE_YMS_NJ001|48|US|1|Advanced Noise Reduction Indicator
0043|GE_YMS_NJ001|49|US|1|Scatter Correction Indicator
0043|GE_YMS_NJ001|4a|DS|3|Recon Center Coordinates
0119|MRSC|1231|IS|1-n|OrthogonalReFormat
0043|GE_YMS_NJ001|50|US|1|Cross-Talk Correction Indicator
0043|GE_YMS_NJ001|51|US|1|Q-Cal Correction Indicator
0043|GE_YMS_NJ001|52|US|1|Afterglow Correction Indicator
0043|GE_YMS_NJ001|53|US|1|Local Decon Correction Indicator
0043|GE_YMS_NJ001|54|DS|1|Scan Start location
0043|GE_YMS_NJ001|55|DS|1|Scan End location
0043|GE_YMS_NJ001|56|IS|1|Detector Row
0043|GE_YMS_NJ001|57|CS|1|Tube Focus
0043|SIEMENS MED NM|03|FL|1-n|View Dependent Y Shift MHR For Detector 1
0045|GEMS_HELIOS_01|0a|FL|1|Minimum DAS value
0045|GEMS_HELIOS_01|18|SS|1|Number of Views 1B
0045|GEMS_HELIOS_01|1a|SS|1|Air Calibration Time
0045|GEMS_HELIOS_01|1b|SS|1|Phantom Calibration Date
0045|GEMS_HELIOS_01|1c|SS|1|Phantom Calibration Time
0045|GEMS_HELIOS_01|1d|SS|1|Z Slope Calibration Date
0045|GEMS_HELIOS_01|1e|SS|1|Z Slope Calibration Time
0045|GEMS_HELIOS_01|1f|SS|1|Cross Talk Calibration Date
0045|GEMS_HELIOS_01|20|SS|1|Cross Talk Calibration Time
0045|GEMS_HELIOS_01|34|CS|1|ActualPctRpeakDelay
0045|GEMS_HELIOS_01|3f|IS|1|RPeakTimeDelay
0045|GEMS_HELIOS_01|44|IS|1|ActualRPeakTimeDelay
0045|GEMS_HELIOS_01|45|ST|1|CardiacScanOption
0049|GEMS_CT_CARDIAC_001|01|SQ|1|CT Cardiac Sequence
0049|GEMS_CT_CARDIAC_001|05|CS|1|MaxHeartRatePriorToConfirm
0049|GEMS_CT_CARDIAC_001|16|SH|1|EkgGatingType
0049|GEMS_CT_CARDIAC_001|1b|FL|1|Ekg Wave Time Off First Data Point
0049|GEMS_CT_CARDIAC_001|22|CS|1|TemporalAlg
0049|GEMS_CT_CARDIAC_001|23|CS|1|PhaseLocation
0049|GEMS_CT_CARDIAC_001|24|OW|1|PreBlendedCycle1
0049|GEMS_CT_CARDIAC_001|25|OW|1|PreBlendedCycle2
0049|GEMS_CT_CARDIAC_001|26|CS|1|CompressionAlg
004b|GEMS_HINO_CT_01|01|DS|1-n|Beam Thickness
004b|GEMS_HINO_CT_01|02|DS|1-n|R Time
004b|GEMS_HINO_CT_01|03|IS|1|HBC number
004b|GE_YMS_NJ001|01|DS|1-n|Beam Thickness
004b|GE_YMS_NJ001|02|DS|1-n|R Time
004b|GE_YMS_NJ001|03|IS|1|HBC number
0051|GEHC_CT_ADVAPP_001|01|SQ|1|CTVESSequence
0051|GEMS_FUNCTOOL_01|01|LO|1|Group Name
0051|GEMS_FUNCTOOL_01|08|SL|1|Color Ramp Index
0053|GEHC_CT_ADVAPP_001|01|FL|1-n|MultiEnergyNoiseRedBlendingFact
0053|GEHC_CT_ADVAPP_001|02|FL|1-n|MultiEnergyNoiseRedScaleFact
0053|GEHC_CT_ADVAPP_001|03|IS|2|MultiEnergyMDTransformEnergies
0053|GEHC_CT_ADVAPP_001|21|IS|1|TableSpeedNotReachesTargetFlag
0053|GEHC_CT_ADVAPP_001|60|SH|1|Recon Flip RotateA nno
0053|GEHC_CT_ADVAPP_001|63|CS|1|Image Position Patient Setting
0053|GEHC_CT_ADVAPP_001|64|IS|1|Shutter Mode
0053|GEHC_CT_ADVAPP_001|65|IS|1|Shutter Mode Percent
0053|GEHC_CT_ADVAPP_001|66|LO|1|Image Browser Annotation
0053|GEHC_CT_ADVAPP_001|67|IS|1|Overlapped Recon Flag
0053|GEHC_CT_ADVAPP_001|68|IS|1|Row Number Anotation Flag
0053|GEHC_CT_ADVAPP_001|70|IS|1|MultiEnergySourceCount
0053|GEHC_CT_ADVAPP_001|71|LO|1|MultiEnergyScanType
0053|GEHC_CT_ADVAPP_001|72|LO|1|MultiEnergyReconType
0053|GEHC_CT_ADVAPP_001|73|LO|1|MultiEnergyImageType
0053|GEHC_CT_ADVAPP_001|74|LO|1|MultiEnergyMaterialType
0053|GEHC_CT_ADVAPP_001|75|DS|1|MonchromaticEnergy
0053|GEHC_CT_ADVAPP_001|76|DS|1|multiEnergyWeightedSubractionWidth1
0053|GEHC_CT_ADVAPP_001|77|DS|1|MultiEnergyWeightedSubractionWidth2
0053|GEHC_CT_ADVAPP_001|78|LO|1|MultiEnergyWeightedSubtractionType
0053|GEHC_CT_ADVAPP_001|79|LO|1|MultiEnergyAcqMethod
0053|GEHC_CT_ADVAPP_001|7a|SH|1|MultiEnergyFeatAnnotName
0053|GEHC_CT_ADVAPP_001|7b|SH|1|MultiEnergyNoiseReduced
0053|GEHC_CT_ADVAPP_001|7c|LO|1|MultiEnergyNoiseReducdeMethod
0053|GEHC_CT_ADVAPP_001|7d|LO|1|SubOptimalIQString
0053|GEHC_CT_ADVAPP_001|7e|DS|1|MultiEnergyHighLowRatio
0053|GEHC_CT_ADVAPP_001|83|DS|1|AnnotationmA
0053|GEHC_CT_ADVAPP_001|84|DS|1|CommandedFirstkVp
0053|GEHC_CT_ADVAPP_001|85|DS|1|CommandedFirstmA
0053|GEHC_CT_ADVAPP_001|86|DS|1|CommandedSecondkVp
0053|GEHC_CT_ADVAPP_001|87|DS|1|CommandedSecondmA
0053|GEHC_CT_ADVAPP_001|88|SH|1|MultiEnergyKVAnnotName
0053|GEHC_CT_ADVAPP_001|89|SH|1|MultiEnergyKVUnitLabel
0053|GEHC_CT_ADVAPP_001|8a|LO|1|MaterialType#1
0053|GEHC_CT_ADVAPP_001|8b|LO|1|MaterialType#2
0053|GEHC_CT_ADVAPP_001|8c|LO|1|GSIScanModePreset
0053|GEHC_CT_ADVAPP_001|8d|IS|1|MonoWindowLow
0053|GEHC_CT_ADVAPP_001|8e|IS|1|MonoWindoHigh
0053|GEHC_CT_ADVAPP_001|8f|FL|1-143|MD1AttenuationCurve
0053|GEHC_CT_ADVAPP_001|92|DS|1|MD1intercept
0053|GEHC_CT_ADVAPP_001|93|DS|1|MD1slope
0053|GEHC_CT_ADVAPP_001|95|OW|1|MD1supportData
0053|GEHC_CT_ADVAPP_001|96|OW|1|MD2supportData
0053|GEHC_CT_ADVAPP_001|97|OW|1|NM1data
0053|GEHC_CT_ADVAPP_001|98|DS|1|MD2intercept
0053|GEHC_CT_ADVAPP_001|99|DS|1|MD2slope
0053|GEHC_CT_ADVAPP_001|9a|OW|1|NM2data
0053|GEHC_CT_ADVAPP_001|9b|FL|1-143|MD2attenuationCurve
0053|GEHC_CT_ADVAPP_001|9c|SH|1|GSIdataVersion
0053|GEHC_CT_ADVAPP_001|9e|IS|1|MultiEnergyNumNoiseRedPair
0053|GEHC_CT_ADVAPP_001|9f|LO|1-n|MultiEnergyNoiseRedPairString
0055|SIEMENS MED NM|04|SS|1|Prompt Window Width
0057|SIEMENS MED NM|01|LO|1|Syngo MI DICOM Original Image Type
0061|SIEMENS MED NM|0f|FL|1-n|X Focal Scaling
0061|SIEMENS MED NM|23|FL|1-n|Recon Selected Angular Range
0061|SIEMENS MED NM|52|LT|1|LowRes CT Series UID
0071|MMCPrivate|01|FL|1|ForegroundTransparency
0071|MMCPrivate|02|LO|1|IsDisplayBackgroundImage
0071|MMCPrivate|03|FL|1|ForegroundHorizontalShift
0071|MMCPrivate|04|FL|1|ForegroundVerticalShift
0119|MRSC|1240|IS|1|LPCCVersion
0071|MMCPrivate|05|FL|1|ForegroundRotationAngle
0071|MMCPrivate|06|FL|1|ForegroundMagnification
0071|MMCPrivate|07|OB|1|ApplicationData
00e1|ELSCINT1|21|DS|1|DLP Total
00e1|ELSCINT1|c2|UI|1|Unknown
0117|MRSC|10|SQ|1|PESERParameterSequence
0117|MRSC|12|CS|1|PESERParameterType
0117|MRSC|14|LO|1|PESERParameterName
0117|MRSC|16|LO|1|PESERParameterDescription
0117|MRSC|18|DS|1-n|PESERParameterFloatingValue
0117|MRSC|19|IS|1-n|PESERParameterIntegerValue
0117|MRSC|1a|LO|1-n|PESERParameterStringValue
0117|MRSC|20|SQ|1|VOISequence
0117|MRSC|22|SQ|1|OmitVOISequence
0117|MRSC|24|SQ|1|ImageQualitySequence
0117|MRSC|30|IS|1|NumberAcquiredTimePoints
0117|MRSC|31|DS|1|AcquisitionDuration
0117|MRSC|32|DS|1-n|AcquisitionStartTimes
0117|MRSC|33|TM|1|InjectionTime
0117|MRSC|34|DS|1-n|EffectiveAcquisitionDelay
0117|MRSC|35|IS|3|SERTimingIndices
0117|MRSC|3a|LO|1|AcquisitionTimingMethod
0117|MRSC|3b|LT|1|AcquisitionTimingComments
0117|MRSC|41|IS|1|ROIVOILPSFlag
0117|MRSC|42|DS|3|VOILPSCenter
0117|MRSC|43|DS|3|VOILPSWidthHalfLength
0117|MRSC|44|DS|3|VOILPSHeightHalfLength
0117|MRSC|45|DS|3|VOILPSDepthHalfLength
0117|MRSC|46|CS|1|VOILPSType
0117|MRSC|50|US|3|ProjectedROINPixels
0117|MRSC|51|IS|1|ProjectedROIProjectionAxis
0117|MRSC|52|IS|1|ProjectedROITransposeFlag
0117|MRSC|53|US|1-n|ProjectedROIXVerts
0117|MRSC|54|US|1-n|ProjectedROIYVerts
0117|MRSC|55|US|2|ProjectedROIZRange
0117|MRSC|56|CS|1|ProjectedROIType
0117|MRSC|5a|LO|1|ProjectedROILabel
0117|MRSC|a1|US|3|FTVPixelLimitsStart
0117|MRSC|a2|US|3|FTVPixelLimitsEnd
0117|MRSC|a3|CS|1|FTVBackgroundMethod
0117|MRSC|a4|DS|1|FTVBackgroundThreshold
0117|MRSC|b0|SQ|1|FTVSequence
0117|MRSC|b1|DS|1|FTVSERMinimum
0117|MRSC|b2|DS|1|FTVSERMaximum
0117|MRSC|b3|IS|1|FTVPixelCount
0117|MRSC|b4|DS|1|FTVcc
0117|MRSC|b5|LO|1|FTVLabel
0117|MRSC|c0|CS|1|QualityControlType
0117|MRSC|c1|LO|1|QualityControlFactor
0117|MRSC|c2|DS|1|QualityControlValue
0117|MRSC|c3|CS|1|QualityControlMeaning
0117|MRSC|c4|LT|1|QualityControlComment
0117|MRSC|c5|CS|1|ProtocolCompliantFlag
0117|MRSC|c6|LO|1-n|ProtocolNotCompliantReasons
0117|MRSC|c7|CS|1|ImagesAnalyzable
0117|MRSC|c8|LO|1-n|ProtocolNotCAnalyzableReasons
0119|MRSC|1000|DS|1|Version
0119|MRSC|1006|DS|1|MinimumPixelValue
0119|MRSC|1007|DS|1|MaximumPixelValue
0119|MRSC|1010|IS|1|PixelDataType
0119|MRSC|1011|IS|1-n|ImageIDNumbers
0119|MRSC|1012|IS|1-n|ParameterDims
0119|MRSC|1013|CS|1-n|VariableParameter
0119|MRSC|1020|LO|1-n|SourceFileNames
0119|MRSC|1021|IS|1|SourceCropFlag
0119|MRSC|1022|IS|6|SourceCropLimits
0119|MRSC|1241|LO|1|LPCCFilename
0119|MRSC|1023|UI|1-n|SourceFileUIDs
0119|MRSC|1024|IS|1-n|SourceVolumeIndices
0119|MRSC|1025|LO|1-n|SourceVolumeLabels
0119|MRSC|1030|DS|9|DirectionCosines
0119|MRSC|1031|CS|3|PatientOrientation3
0119|MRSC|1041|DS|1-n|SlicePosition
0119|MRSC|1050|LO|1-n|VolumeLabels
0119|MRSC|1051|DA|1-n|AcquisitionDate
0119|MRSC|1060|LO|1|SecCptrUser
0119|MRSC|1061|LO|1|SecCptrApplication
0119|MRSC|1070|AT|1-n|VariableParamTags
0119|MRSC|1071|CS|1-n|VariableParamNames
0119|MRSC|1080|DS|1-n|TR
0119|MRSC|1081|DS|1-n|TE
0119|MRSC|10a0|DS|1-n|DIFF_GRAD_X
0119|MRSC|10a1|DS|1-n|DIFF_GRAD_Y
0119|MRSC|10a2|DS|1-n|DIFF_GRAD_Z
0119|MRSC|10a3|DS|1-n|DIFF_PW_X
0119|MRSC|10a4|DS|1-n|DIFF_PW_Y
0119|MRSC|10a5|DS|1-n|DIFF_PW_Z
0119|MRSC|10a6|DS|1-n|DIFF_TIME_X
0119|MRSC|10a7|DS|1-n|DIFF_TIME_Y
0119|MRSC|10a8|DS|1-n|DIFF_TIME_Z
0119|MRSC|10a9|DS|1-n|DiffBValues
0119|MRSC|10b0|LO|1|CoilCorrectionMethod
0119|MRSC|10b1|IS|1|PolyFitOrder
0119|MRSC|10b2|DS|1-n|PolyFitCoeff
0119|MRSC|1100|DS|1|FitMapModuleVersion
0119|MRSC|1101|LO|1-n|SourceFileNames
0119|MRSC|1102|IS|1-n|SourceVolumeIndices
0119|MRSC|1103|DS|1-n|ParameterValues
0119|MRSC|1104|AT|1|ParameterTag
0119|MRSC|1105|UI|1-n|SourceFileUIDs
0119|MRSC|1106|LO|1-n|SourceFileDirectory
0119|MRSC|1107|IS|1|SourceDataInPlaceFlag
0119|MRSC|1108|IS|1-n|ResultVolumeindices
0119|MRSC|1109|IS|1|SMOOTHBoxcarAverageKernel
0119|MRSC|110c|LO|1|FitICFunction
0119|MRSC|110d|LO|1|FitFormulaProcedure
0119|MRSC|110e|LO|1|FittingProgram
0119|MRSC|110f|IS|1|FittingProgramVersion
0119|MRSC|1110|CS|1|FitType
0119|MRSC|1111|IS|1|SetICFlag
0119|MRSC|1112|DS|1-n|InitialConditions
0119|MRSC|1113|DS|1-n|FitMapScaleFactors
0119|MRSC|1120|IS|1|ThresholdingFlag
0119|MRSC|1121|DS|1|Threshold
0119|MRSC|1122|IS|1|MaskCompression
0119|MRSC|1123|OB|1-n|FitMapMask
0119|MRSC|1124|OB|1-n|FitMapPntThreshMap
0119|MRSC|1125|ST|1|PixelMaskCheckString
0119|MRSC|1250|IS|1|LPCCFilter_type
0119|MRSC|1251|DS|1|LPCCMean_Multiplier
0119|MRSC|1260|DS|1|SACoilCorrectionIncrement
0119|MRSC|1261|IS|1|SACoilCorrectionVersion
0119|MRSC|1270|DS|1|SACoilCorrectionParams_Angle_deg
0119|MRSC|1271|DS|1|SACoilCorrectionParams_Offset_in
0119|MRSC|12a0|LO|1|MinVarFiltSid
0119|MRSC|12a1|LO|1|MinVarFiltPath
0119|MRSC|12a2|IS|1|MinVarFiltMax_images
0119|MRSC|12a3|IS|2|MinVarFiltId_locs
0119|MRSC|12a4|LO|1|MinVarFiltScript_name
0119|MRSC|12a5|IS|1|MinVarFiltSave_masks
0119|MRSC|12a6|IS|1|MinVarFiltSave_idf
0119|MRSC|12a7|LO|1|MinVarFiltMask
0119|MRSC|12a8|LO|1|MinVarFiltIdfmask
0119|MRSC|12a9|LO|1|MinVarFiltImage
0119|MRSC|12b0|IS|1|MinVarFiltOutput_type
0119|MRSC|12b1|IS|1|MinVarFiltOutput_ftype
0119|MRSC|12b2|LO|1|MinVarFiltScaling
0119|MRSC|14|UI|1|SERMaskFileUID
0119|MRSC|1400|LO|1|MIPsSid
0119|MRSC|1401|UI|1|MIPsUID
0119|MRSC|1402|TM|1|MIPsTime
0119|MRSC|1403|DA|1|MIPsDate
0119|MRSC|1404|IS|1|MIPsVersion
0119|MRSC|1405|IS|1|MIPsVolume
0119|MRSC|1406|IS|1|MIPsOrtho
0119|MRSC|1407|IS|1|MIPsMaskedFlag
0119|MRSC|1408|IS|1|MIPsSubtractVolume
0119|MRSC|1410|UL|1-n|MIPsProtectPixels
0119|MRSC|1411|UL|1-n|MIPsIgnorePixels
0119|MRSC|1412|IS|1|MIPsProjectFlag
0119|MRSC|1413|IS|1-n|MIPsProjectPlaneIndices
0119|MRSC|1500|LO|1|SERSid
0119|MRSC|1501|UI|1|SERUID
0119|MRSC|1503|DA|1|SERDate
0119|MRSC|1504|IS|1|SERVersion
0119|MRSC|1505|IS|3|SERTimePoints
0119|MRSC|1506|IS|1|SERByteScaled
0119|MRSC|1507|DS|1|SERBackground
0119|MRSC|1508|DS|1|SERThreshold
0119|MRSC|1509|DS|1|SERMaximum
0119|MRSC|150a|IS|1|SERMinConPixels
0119|MRSC|150b|IS|1|SERCorrectFlag
0119|MRSC|150c|DS|2|SERAcqTimes
0119|MRSC|150d|DS|2|SERTargetTimes
0119|MRSC|150e|DS|1|SERTimeTolerance
0119|MRSC|150f|DS|4|SERCorrectionParams
0119|MRSC|1510|LO|1|SERImageType
0119|MRSC|1511|IS|1-n|SEROffsets
0119|MRSC|1512|LO|1|SERMaskFileName
0119|MRSC|1513|DS|1|SERMaskChecksum
0119|MRSC|18|IS|3|GAINS
0119|MRSC|27|IS|1-n|ByteScaleMinMaxTop
0119|MRSC|28|IS|1-n|GlobalThreshold
0119|MRSC|29|DS|1-n|IntensityScale
0119|MRSC|32|IS|1-n|REBIN
0119|MRSC|33|DS|1-n|WhiteTopHat
0119|MRSC|34|IS|1-n|HistEqual
0119|MRSC|35|IS|1-n|Crop
0119|MRSC|36|DS|1-n|LPCoil
0119|MRSC|38|DS|3|PixelGap
0119|MRSC|42|DS|1-n|LPCCBandwidth
0119|MRSC|43|DS|1|LPCCNoise_factor
0119|MRSC|44|DS|1|LPCCNoise_level
0119|MRSC|45|IS|1|LPCCNoise_mode
0119|MRSC|46|IS|1|LPCCDirection
0119|MRSC|47|IS|1|LPCCEdge_fill
0119|MRSC|48|IS|1|LPCCMean_fill
0119|MRSC|49|IS|1|LPCCPixelsearch
0119|MRSC|4a|DS|1|LPCCIntensity_scale
0119|MRSC|4b|IS|1|LPCCThreed
0119|MRSC|4c|LO|1|LPCCRoi_mask
0119|MRSC|4d|IS|2|LPCCMask_slices
0119|MRSC|4e|IS|1|LPCCSlice_pad
0119|MRSC|4f|IS|1|LPCCSave_type
0119|MRSC|52|TM|1-n|AcquisitionTime
0119|MRSC|62|DA|1|SACoilCorrectionCorr_date
0119|MRSC|63|TM|1|SACoilCorrectionCorr_time
0119|MRSC|64|LO|1|SACoilCorrectionMethod
0119|MRSC|65|DS|1-n|SACoilCorrectionOrigin
0119|MRSC|66|DS|1-n|SACoilCorrectionAxis_cos
0119|MRSC|67|IS|1|SACoilCorrectionNumber
0119|MRSC|68|LO|1|SACoilCorrectionSid
0119|MRSC|69|DS|1-n|SACoilCorrectionRange
0119|MRSC|6a|FD|1-n|SACoilCorrectionSa_value
0119|MRSC|6b|IS|1|SACoilCorrectionAxis_flag
0119|MRSC|6c|IS|1-n|SACoilCorrectionSample_number
0119|MRSC|6d|LO|1|SACoilCorrectionParams_SID
0119|MRSC|6e|IS|1|SACoilCorrectionParams_Version
0119|MRSC|6f|DS|1|SACoilCorrectionParams_Rot_axis_off
0119|MRSC|72|DS|1-n|SACoilCorrectionParams_Plane_cos_ref
0119|MRSC|73|DS|1-n|SACoilCorrectionParams_Lps_ref
0119|MRSC|74|IS|1|SACoilCorrectionParams_Order
0119|MRSC|75|DS|1-n|SACoilCorrectionParams_Coeff
0119|MRSC|76|DA|1|SACoilCorrectionParams_Coeff_date
0119|MRSC|77|LO|1|SACoilCorrectionParams_Coeff_src
0119|MRSC|82|DS|1-n|TI
0119|MRSC|83|DS|1-n|TSL
0119|MRSC|88|DS|1-n|FlipAngle
0119|MRSC|90|DS|1-n|TemporalIndex
0119|MRSC|91|DS|1-n|TemporalValue
0119|MRSC|aa|LO|1-n|MinVarFiltIdfimages
0119|MRSC|ab|LO|1|MinVarFiltOutput_file
0119|MRSC|ac|IS|1|MinVarFiltNum_loops
0119|MRSC|ad|IS|3|MinVarFiltKernel
0119|MRSC|ae|IS|1|MinVarFiltLimit_sliceFlag
0119|MRSC|af|SS|2|MinVarFiltSlice_limits
0119|MRSC|b3|LO|1|MinVarFiltScript
0119|MRSC|b4|LO|1|MinVarFiltLog
0119|MRSC|c0|SQ|1|QCMinimumLimits
0119|MRSC|c1|SQ|1|QCMaximumLimits
0119|MRSC|d0|ST|1|CheckString
0119|MRSC|d1|LO|1-n|Source
0119|MRSC|f0|OB|1-n|SampleHeader
0119|MRSC|ff|DS|1-n|UserInfo
01e1|ELSCINT1|c2|UI|1|GT Gating UID
1001|BrainWave: 1.2.840.113819.3|11|SH|1|DICOM Implementation Version
2001|BrainWave: 1.2.840.113819.3|10|UI|1|DICOM Implementation UID
2001|BrainWave: 1.2.840.113819.3|12|UI|1|Within-DICOM-Implementation SOP Instance UID
2001|BrainWave: 1.2.840.113819.3|13|SH|1|Application Name
2001|BrainWave: 1.2.840.113819.3|14|SH|1|Application Version
2001|BrainWave: 1.2.840.113819.3|15|SH|1|Compatibility Version
2001|BrainWave: 1.2.840.113819.3|21|UI|1-n|Referenced Series UID
2001|BrainWave: 1.2.840.113819.3|31|US|1|Number of Objects Averaged
2001|BrainWave: 1.2.840.113819.3|41|US|1|Number of Expected Time Points
2001|BrainWave: 1.2.840.113819.3|51|US|1|Number of Slices Per Volume
2001|BrainWave: 1.2.840.113819.3|60|US|1|BW Image Type
2001|BrainWave: 1.2.840.113819.3|61|US|1|Experiment Type
2001|BrainWave: 1.2.840.113819.3|71|UI|1|Paradigm UID
2001|BrainWave: 1.2.840.113819.3|72|LO|1|Paradigm Name
2001|BrainWave: 1.2.840.113819.3|73|ST|1|Paradigm Description
2001|BrainWave: 1.2.840.113819.3|80|OB|1|Contrast
2001|BrainWave: 1.2.840.113819.3|81|FL|1-n|Regressor Values
2001|BrainWave: 1.2.840.113819.3|86|US|1|Number of Degrees of Freedom
2001|BrainWave: 1.2.840.113819.3|8a|FL|1|Z Threshold
2001|BrainWave: 1.2.840.113819.3|8b|FL|1|p Threshold
2001|BrainWave: 1.2.840.113819.3|90|OB|1|Processing Parameters
2001|BrainWave: 1.2.840.113819.3|91|OB|1|Motion Plot
2001|BrainWave: 1.2.840.113819.3|92|OB|1|ROIs
2001|BrainWave: 1.2.840.113819.3|93|OB|1|Tracts
2001|BrainWave: 1.2.840.113819.3|94|OB|1|Report
2001|BrainWave: 1.2.840.113819.3|95|OB|1|Response Data
2001|BrainWave: 1.2.840.113819.3|a0|FL|1-n|Motion Parameters
2001|BrainWave: 1.2.840.113819.3|a1|FL|1-n|Registration Parameters
2001|BrainWave: 1.2.840.113819.3|a2|FL|1-n|Subject Data
2001|BrainWave: 1.2.840.113819.3|b0|OB|1|DTI Parameters
2001|BrainWave: 1.2.840.113819.3|c0|OB|1|Paradigm Info
2001|Philips Imaging DD 001|01|FL|1|ChemicalShift
2001|Philips Imaging DD 001|02|IS|1|ChemicalShiftNumberMR
2001|Philips Imaging DD 001|03|FL|1|DiffusionB-Factor
2001|Philips Imaging DD 001|04|CS|1|DiffusionDirection
2001|Philips Imaging DD 001|06|CS|1|ImageEnhanced
2001|Philips Imaging DD 001|07|CS|1|ImageTypeEDES
2001|Philips Imaging DD 001|08|IS|1|PhaseNumber
2001|Philips Imaging DD 001|09|FL|1|Image Prepulse Delay
2001|Philips Imaging DD 001|0a|IS|1|SliceNumberMR
2001|Philips Imaging DD 001|0b|CS|1|SliceOrientation
2001|Philips Imaging DD 001|0c|CS|1|Arrhythmia Rejection
2001|Philips Imaging DD 001|0e|CS|1|Cardiac Cycled
2001|Philips Imaging DD 001|0f|SS|1|Cardiac Gate Width
2001|Philips Imaging DD 001|10|CS|1|Cardiac Sync
2001|Philips Imaging DD 001|11|FL|1|DiffusionEchoTime
2001|Philips Imaging DD 001|12|CS|1|DynamicSeries
2001|Philips Imaging DD 001|13|SL|1|EPIFactor
2001|Philips Imaging DD 001|14|SL|1|NumberOfEchoes
2001|Philips Imaging DD 001|15|SS|1|NumberOfLocations
2001|Philips Imaging DD 001|16|SS|1|NumberOfPCDirections
2001|Philips Imaging DD 001|19|CS|1|PartialMatrixScanned
2001|Philips Imaging DD 001|1b|FL|1|PrepulseDelay
2001|Philips Imaging DD 001|1c|CS|1|PrepulseType
2001|Philips Imaging DD 001|1d|IS|1|ReconstructionNumberMR
2001|Philips Imaging DD 001|1f|CS|1|RespirationSync
2001|Philips Imaging DD 001|21|CS|1|SPIR
2001|Philips Imaging DD 001|22|FL|1|WaterFatShift
2001|Philips Imaging DD 001|23|DS|1|FlipAnglePhilips
2001|Philips Imaging DD 001|25|SH|1|EchoTimeDisplayMR
2001|Philips Imaging DD 001|2d|SS|1|StackNumberOfSlices
2001|Philips Imaging DD 001|32|FL|1|StackRadialAngle
2001|Philips Imaging DD 001|33|CS|1|StackRadialAxis
2001|Philips Imaging DD 001|35|SS|1|StackSliceNumber
2001|Philips Imaging DD 001|36|CS|1|StackType
2001|Philips Imaging DD 001|58|UL|1|Contrast Transfer Taste
2001|Philips Imaging DD 001|5f|SQ|1-n|StackSequence
2001|Philips Imaging DD 001|60|SL|1|NumberOfStacks
2001|Philips Imaging DD 001|61|CS|1|SeriesTransmitted
2001|Philips Imaging DD 001|63|CS|1|ExaminationSource
2001|Philips Imaging DD 001|7b|IS|1|AcquisitionNumber
2001|Philips Imaging DD 001|81|IS|1|NumberOfDynamicScans
2001|Philips Imaging DD 001|a1|CS|1|Is Raw Image
2001|Philips Imaging DD 001|c8|LO|1|Exam Card Name
2001|Philips Imaging DD 001|f1|FL|6|Prospective Motion Correction
2001|Philips Imaging DD 001|f2|FL|6|Retrospective Motion Correction
2005|Philips MR Imaging DD 001|20|SL|1|NumberOfChemicalShifts
2005|Philips MR Imaging DD 001|a1|CS|1|SyncraScanType
2005|Philips MR Imaging DD 001|b0|FL|1|Diffusion Direction RL
2005|Philips MR Imaging DD 001|b1|FL|1|Diffusion Direction AP
2005|Philips MR Imaging DD 001|b2|FL|1|Diffusion Direction FH
50f1|FDMS 1.0|06|CS|1|Energy Subtraction Parameter
50f1|FDMS 1.0|07|CS|1|Subtraction Registration Result
50f1|FDMS 1.0|08|CS|1|Energy Subtraction Parameter 2
50f1|FDMS 1.0|09|SL|1|Afin Conversion Coefficient
50f1|FDMS 1.0|20|CS|1|Image Processing Modification Flag
7001|GEMS_MR_RAW_01|01|OB|1|rdb_hdr_rec
7001|GEMS_MR_RAW_01|02|OB|1|rdb_hdr_per_pass_tab
7001|GEMS_MR_RAW_01|03|OB|1|rdr_hdr_unlock_raw
7001|GEMS_MR_RAW_01|04|OB|1|rdb_hdr_data_acq_tab
7001|GEMS_MR_RAW_01|05|OB|1|rdb_hdr_nex_tab
7001|GEMS_MR_RAW_01|06|OB|1|rdb_hdr_nex_abort_tab
7001|GEMS_MR_RAW_01|07|OB|1|rdb_hdr_tool
7001|GEMS_MR_RAW_01|08|OB|1|rdb_raw_data
7001|GEMS_MR_RAW_01|09|OB|1|SSP save
7001|GEMS_MR_RAW_01|0a|OB|1|UDA save
7001|GEMS_MR_RAW_01|0b|OB|1|rdb_chemsat_data
7005|TOSHIBA_MEC_CT3|00|OB|1|CT Private Data 1
7005|TOSHIBA_MEC_CT3|03|SH|1|Cardiac R-R Mean Time
7005|TOSHIBA_MEC_CT3|04|SH|1|Cardiac Reconstruction Getting Phase in Percent
7005|TOSHIBA_MEC_CT3|05|SH|1|Cardiac Reconstruction Getting Phase in ms
7005|TOSHIBA_MEC_CT3|06|SH|1|Cardiac Reconstruction Mode
7005|TOSHIBA_MEC_CT3|07|DS|1-n|Reconstruction Center
7005|TOSHIBA_MEC_CT3|08|DS|1|Detector Slice Thickness in mm
7005|TOSHIBA_MEC_CT3|09|LO|1|Number of Detector rows to Reconstruct
7005|TOSHIBA_MEC_CT3|0a|DS|1|Table Speed in mm/rot
7005|TOSHIBA_MEC_CT3|0b|SH|1|Filter
7005|TOSHIBA_MEC_CT3|0c|SH|1|Reconstruction Correction Type
7005|TOSHIBA_MEC_CT3|0d|SH|1|Organ
7005|TOSHIBA_MEC_CT3|0e|SH|1|File Type Remarks
7005|TOSHIBA_MEC_CT3|0f|SH|1|Direction (head or feet first)
7005|TOSHIBA_MEC_CT3|10|OB|1|CT Private Data 2
7005|TOSHIBA_MEC_CT3|11|LT|1|Series Comment
7005|TOSHIBA_MEC_CT3|12|SH|1|Position (supine or prone)
7005|TOSHIBA_MEC_CT3|13|US|1|Expert Plan Number
7005|TOSHIBA_MEC_CT3|14|US|1|Reconstruction ROI Number
7005|TOSHIBA_MEC_CT3|15|US|1|Special Helical Acquisition Number
7005|TOSHIBA_MEC_CT3|16|UI|1|Volume UID
7005|TOSHIBA_MEC_CT3|17|US|1|Total Frame Count in the Volume
7005|TOSHIBA_MEC_CT3|18|US|1|Frame Number
7005|TOSHIBA_MEC_CT3|19|UL|1|Frame Sort Key
7005|TOSHIBA_MEC_CT3|1a|US|1|Frame Sort Order
7005|TOSHIBA_MEC_CT3|1b|SH|1|Convolution Kernel for Series Record
7005|TOSHIBA_MEC_CT3|1c|LO|1|Contrast/Bolus Agent for Series Record
7005|TOSHIBA_MEC_CT3|1d|UL|1|Reconstruction Number
7005|TOSHIBA_MEC_CT3|1e|UL|1|Raw Data Number
7005|TOSHIBA_MEC_CT3|1f|LO|1|Volume Number
7005|TOSHIBA_MEC_CT3|20|UL|1|Local Series Number
7005|TOSHIBA_MEC_CT3|21|LO|1|Decrease in Artifact Filter
7005|TOSHIBA_MEC_CT3|22|DS|1|Reconstruction Interval
7005|TOSHIBA_MEC_CT3|23|DS|1|Pitch Factor
7005|TOSHIBA_MEC_CT3|24|DA|1|AcquisitionDateOfNRA
7005|TOSHIBA_MEC_CT3|25|UL|1|Large Data File Attribute
7005|TOSHIBA_MEC_CT3|26|CS|40915|Large Data File Name
7005|TOSHIBA_MEC_CT3|28|SQ|1|Enhanced CT Private Sequence
7005|TOSHIBA_MEC_CT3|29|UI|1|Frame UID
7005|TOSHIBA_MEC_CT3|30|CS|1|Main Modality in Study
7005|TOSHIBA_MEC_CT3|35|DS|2|Scan Range
7005|TOSHIBA_MEC_CT3|36|OB|1|CT Private Data 3
7005|TOSHIBA_MEC_CT3|37|IS|1|Total Frames
7005|TOSHIBA_MEC_CT3|38|IS|1|Start Frame
7005|TOSHIBA_MEC_CT3|39|IS|1|End Frame
7005|TOSHIBA_MEC_CT3|40|FD|1|DLP
7005|TOSHIBA_MEC_CT3|41|SH|1|Row Slice Information
7005|TOSHIBA_MEC_CT3|42|US|1|Local Frame Number
7005|TOSHIBA_MEC_CT3|43|DS|3|Volume Vector
7005|TOSHIBA_MEC_CT3|44|US|1|Volume Type
7005|TOSHIBA_MEC_CT3|45|DS|1|Relative Table Position of 4D Volume
7005|TOSHIBA_MEC_CT3|46|DS|1|Absolute Table Position of 4D Volume
7005|TOSHIBA_MEC_CT3|47|DS|1|Slice Pitch of 4D Volume
7005|TOSHIBA_MEC_CT3|48|LO|1|Respiratory Gating Information
7005|TOSHIBA_MEC_CT3|49|SH|1|Respiratory Phase
7005|TOSHIBA_MEC_CT3|f1|CS|1|Protect Mark for Image, Curve or Private Record
7005|TOSHIBA_MEC_CT3|f2|CS|1|Protect Mark for Series Record
7005|TOSHIBA_MEC_CT3|f3|CS|1|Protect Mark for Study Record
700d|TOSHIBA_MEC_MR3|00|DS|1|Scale Factor
700d|TOSHIBA_MEC_MR3|01|OB|1|Acquisition Order
700d|TOSHIBA_MEC_MR3|02|DS|1|Orientation Vector
700d|TOSHIBA_MEC_MR3|03|SS|1|Flip Flag
700d|TOSHIBA_MEC_MR3|04|OB|1|Rotate Information
700d|TOSHIBA_MEC_MR3|05|DS|1|FOV
700d|TOSHIBA_MEC_MR3|06|US|1|Image Matrix
700d|TOSHIBA_MEC_MR3|07|OB|1|Image Information
700d|TOSHIBA_MEC_MR3|08|OB|1|Original Data
700d|TOSHIBA_MEC_MR3|09|SS|1|Original Data Flag
700d|TOSHIBA_MEC_MR3|80|US|N|Number of PAC channel
700d|TOSHIBA_MEC_MR3|81|US|N|Reference mode
700d|TOSHIBA_MEC_MR3|82|SQ|N|Gain value group for MRS
700d|TOSHIBA_MEC_MR3|88|UL|N|Flag of water Sat pulse
700d|TOSHIBA_MEC_MR3|89|FL|N|Selected contrast TE
700d|TOSHIBA_MEC_MR3|8a|SQ|N|Raw Data Set Sequence
700d|TOSHIBA_MEC_MR3|91|FL|N|Receiver gain of prescan
7053|Philips PET Private Group|00|DS|1|SUV Factor
7053|Philips PET Private Group|01|OB|1|Private Data
7053|Philips PET Private Group|02|OB|1|Private Data
7053|Philips PET Private Group|03|ST|1|Original File Name
7053|Philips PET Private Group|05|LO|1|Worklist Info File Name
7053|Philips PET Private Group|06|OB|1|Unknown
7053|Philips PET Private Group|07|SQ|1|Unknown
7053|Philips PET Private Group|09|DS|1|Activity Concentration Scale Factor
7053|Philips PET Private Group|13|SS|1|Unknown
7053|Philips PET Private Group|14|SS|1|Unknown
7053|Philips PET Private Group|15|SS|1|Unknown
7053|Philips PET Private Group|16|SS|1|Unknown
7053|Philips PET Private Group|17|SS|1|Unknown
7053|Philips PET Private Group|18|SS|1|Unknown
7053|Philips PET Private Group|c2|UI|1|Unknown
7fe1|SIEMENS CSA NON-IMAGE|10|OB|1|CSA Data
7fe3|SIEMENS MED NM|14|OW|1|Minimum Pixel in Frame
7fe3|SIEMENS MED NM|15|OW|1|Maximum Pixel in Frame
7fe3|SIEMENS MED NM|29|OW|1|Number of R-Waves in Frame
